<svg xmlns="http://www.w3.org/2000/svg" version="1.1" xmlns:xlink="http://www.w3.org/1999/xlink" width="384" height="384"><svg xmlns="http://www.w3.org/2000/svg" version="1.1" xmlns:xlink="http://www.w3.org/1999/xlink" width="384" height="384" viewBox="0 0 384 384"><image width="384" height="384" xlink:href="data:image/png;base64,iVBORw0KGgoAAAANSUhEUgAAAgAAAAIACAYAAAD0eNT6AAABdGVYSWZNTQAqAAAACAAEAQAABAAAAAEAAAAAAQEABAAAAAEAAAAAh2kABAAAAAEAAAA+ARIABAAAAAEAAAAAAAAAAAACkoYAAgAAARgAAABckggABAAAAAEAAAAAAAAAAHsicmVtaXhfZGF0YSI6W10sInNvdXJjZV90YWdzIjpbXSwidG90YWxfZHJhd190aW1lIjowLCJ0b3RhbF9kcmF3X2FjdGlvbnMiOjAsImxheWVyc191c2VkIjowLCJicnVzaGVzX3VzZWQiOjAsInBob3Rvc19hZGRlZCI6MCwidG90YWxfZWRpdG9yX2FjdGlvbnMiOnt9LCJ0b29sc191c2VkIjp7ImVmZmVjdHMiOjEsInNxdWFyZV9maXQiOjF9LCJpc19zdGlja2VyIjpmYWxzZSwiZWRpdGVkX3NpbmNlX2xhc3Rfc3RpY2tlcl9zYXZlIjp0cnVlLCJjb250YWluc0ZURVN0aWNrZXIiOmZhbHNlfQCYUXLVAAAAAXNSR0IArs4c6QAAAARzQklUCAgICHwIZIgAACAASURBVHic7L33kxxHluf5fe4RkVqUVlAFFEQVNAESJJvN7m0xYq/P5lbdT2d2/92Z3S93P+yenZ3N3szu2fZON5vTFCBAkITWqnTqCPd3P7hHZGShQIKgwjTex6yqsiIj3SMzPP09f8oBQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRAEQRCE50I/9QUIgpDxbb6P/INdhSAIrwWiAAjCjw8BCDA/H473ykFS7gVVW1bGGPXCDRBlCoBSiofHh4+3ANT9421qMeXO+8b2821uvtjrmK2bT5qjx+vWfu08Y60loLHLM5sA3PsAANpWTKSYaJODIDBPnjwxABL/IwqRIHxLRAEQhB8XDaBaqNVmmvXxPVFYniJSdaigqAgBq4CU/17SM0JtKPRBYFhiCwDWMsEyANjsHANLlhU0AxbWWkbangUIxAaGgVSZUO4JB/vH7nmbUzZyZz2rrTAZ/4QGYPzREIqQm2uYVfZYZ29MERRnx60ldi0Qx4hBZK21ZIk5YU4GMNyKYda32psP+pubTwG0cl0KgvACiAIgCD8e5ampqQUKK8cHA3smjMJlReF+rfW4UkGZCQEoGJGWBN51ZcsgBhMYzGBmgIf/ux9YWG8RYGa2DBAT4FtMz0PWEzGnst0/wel1MNhpAwoEC2YaPgfKnclgAgEKRKOKAqVKTfqYiNIrAjGB3JNMBMWWGYCFATOTZVg2TGzZcmwZXct20zLuw/KVYrFwpRzgq2vXPr8LZzYQa4AgvACiAAjCDw8BqNTGF06WiqXfgsLf9mI+bI0tWeZQEWlFDkCNSi8nFN0PI5WSeXYRdu58ZgYRkElrBsgCVvEz7RAAsgRWnDVIdrQ/RirsAVIWqS1AWZ326I4pAqy3Dyh/DARlKNdC1ov7IfbXBZBVYFgwGKwApyO4xb1lzZY1G7AhqKRYUO1KIbylgQ/a2+v/hWz3j0+fPn0KIP7aOyIIgigAgvADQwAqY1NzZ6Pi+L8xRv2iH9uDsTFVpVgRGFqBtNIgRUhiRpIYMBgq0AgiDUUMIgvi3KqbRztIhXOeVCBzJnfdmUzPKhKUa4lTZSH3THae75ez9T1Bsfb9OaWAVd55MRT0yuZViB29k++XCGnTDAanx33rSaKQGIJhMFsFAplIq04UqMcB8GUhTP5j33b+/tHt23cBDHa5H4IgeIKf+gIE4S+ccrM5tVSIxv4utvq3vcQeiq0pKA2qVEsolQJUyyXUqhUQNB4+WMXGxiYsGzTHq5ien0QUKKcEwIL8qnvoUHe2cyYL4h1eeWK/knYvICIQfUOcYdow7/I/jSoe7E+g1JOfKgBEzolAo+3QixjmR16T2hUYTARjgXZ7gFa7j1ZnQK2tHvq9JOjHXE8SlKNATxbL1WrJhv25ubl/fPDgwR3kAhsEQRhFFABB+OEI6vWpubBQ+1tj9V/3Y3twYOKiChnjE1UsLy9iYWEa09PjGKs3kQwY//if/zuuXe2iWA5x6uwxnD13CqVIO5M7Dc3uowqAApMBscaIxKbUnG8BIigQSFEmXzldqOcX+Zm5IA8/I71p5JH2DeVN+7nXfq1LXj33PKbhMSKCSQitVgdra1t4+HgDX315C3duP0Zrs4d4wIExtl4cRBea9dpmqRRuPnjwYANpKoEgCM8gCoAg/GDUGkEhOgsV/vte3xwYGFPUIWNqpoHzby3jl798E4cP78f42BgCCvDo/io+/OBPqNU1lg7vwd/+7Tt48+2zCDWBYLxTPhWKlDPRE5xi8LzV/dBDDyL3iNwRm5rd4QP5mHZpx2YKwG4G/KECkO/S9edcBc9XABQrWBAU3HmWXNjAqEuDnZuBCXGcoN3u48nqJj79+Ap+/9/+jCuf38GTR9sY9I3aanUKtWrpvSAs3108cuTejS+//BBiBRCEXREFQBB+GMKJifISqPCLONZHEmOLiiwmJ+t4680V/Lt//zc4tDSPaq2IgDTWV1v48uoV3L13HfVGASdOH8aJE4dQr2sv/HOCmSzAaocf/5tN+zzy2CsFxIBSXhADBBd1Z/Mi2CsdBIZiwI7kJ6ZKw/AKfGqiN92rnNKw06+QKgAMZ58ALLFPXPSqDXuFxbsZilxAtVrE5EQNC7NTmJmawP9b+SP++MFl3H+4BmM0Hj3dqk2NlX7WbE7frtUeXN/e3n76zbdLEF4/RAEQhO8fqlarTYqqZ5ijtwcDLjEMlUqalg7N4d23T2H56D5UagG0JvR7Ce7ff4jf//6f0Gpt4ujZszh+bAnjkzUobcBInA99ZNX/Tab1nVdETkBTPnmPXJCdtwu4I86SkIpdgOBqDrkVukoDCDNPgxPywNA4oRQxkcosDd7WkCUdcnbpBEVZmqBTMAi+j+wKwcPyACB2JQsCpTA+VsHZsysY9CxarS7WNzfQawNxnOj+wO7vdc2F6em5T7e3t/8BQP/FPyxBeD0QBUAQvn+CsFQ7llh6y1heSqxVQcCYnmngxIlDOHnyEBrNAoAEzMDG+ha++uI6Ln/2Oer1Ok4cP4LFg3tQKBCYEjCMl9sKIyv9TJKmioDKCfhRmG1m6qfcOWny/UjoAHkVgHOCfkfmQN6aQKmA9lKb4YR4mnto4UoOjMYXUibkhzmKnF2+8mdSlo0wzCBgMIgIQQBMTtZx+sxhPHm6irv37uP6tXUMBqBWd1DVIZ2Ympz9m/H19sW1tXsP4SoGCoLgeeHSo4IgvDA1S9EFY+ncILFVC4MgZBxc2oMTpw5jbs8EQK567WBgcPvWA3z80UVsrm9iZeUYjq4cxsRUA6Bh1P9zM3aZ/Mr7mzN62dcM+uYfC7BPO8zqCj3/fF93yP+1ILZZG+nfPCq1JHgNQBGB/P/Dlb9b/TsNwMcgUKokpEGJBlonmJlr4vTZwzh//jiq1QKUYnT7fd3pDOZ6A7zfnKidaTT21V7yXgrCXyyiAAjC94uujY8ftSq8YKEWmUkFITA+UcGJUwdx+MhelMoB0np662tbuPTZFXz26WVUKjWcf/Mc9h6YR6EUgvyKWJOGggY983V1TgEFDQWFryvr4VIA/Vr664Q/LCwMLBtY2G8Q+gxYhvXHLPvX5n44l7WQ5Re4aj94sdi8vBJgXYSgVwJIAUQGUYGx78AM3vvFOcwvjKFQIrC16Hbi0urTrf2N2sTvphbG5iEWT0EYQRQAQfj+UABqhaj6V8zqeGK5DDIoVyOcPnMEp04dwczsGJS2YFjEA4uvvryOzy5eQqfXwclTKzi2chCNZgVQLxa4/rVRALzj51vDWbDgtzvv23T8on3sIFcjgMig0Szi2LFFnHvjKMbGKlCKkSSG4hjlsFD9dUEXTlers2PfrhNB+MtGFABB+P6o1OsTRwY2eNckdo6tVVGkMDFWwRvnT2Df4qxf/ROMIayvt3Dx4hXcvnMX07OT+OVv3sPUTBNBkdy2OsR4keh+Qy4yfzcU+0XzS70dC1eC95uE827npSv8l3ltSpr5sLPAUVol0AJkADIIQ0JzrIx3fnYOB/bPolopgkhRv2+CBw83FhKD9/funT6EbP8hQRBEARCE7wc9ObkwV6k1fg0Kl4yhMoGpXivh2NFFHFs5iPHxGkgB1jL6PYOrX93Glc+vo9vt48ChfTh+8ggq1QhuJ14eutWfJ0Npl5/nnPateYF2v9V5L8qI8eAF3xwxQAZRgbCysoiTK4cwPdkAwSJOEtpudQuKogtBUDlVq9XECiAIHlEABOH7oQqoY5bC37HVUyAEUagwNzuOn/3sHPbtnUGpFIEAmBjYXGvjww8u4u6th5iYmMDpMycwMzuOMFQuKA7Ad7DdZ3wnD8CPxm7C/dljWfzBrlhobTE9Xce58ytYPDCPUjEAwBQnltpdc7iX4MLCwv4jz+lQEF47RAEQhO+OHpuZ2WfC8O1+gpODxJSImMYmqlhePoA33zqJsWYZgQJgCb12jFvX7+HTjy/DGIsTx1dw/o3TKBY0NAE6jZBHmn//khDAym/M96OKPF8eGBrfPMXsdnEabn+BFwtqzBwFxNChwdHlAzhx8hDm5iYQaGdxWd9sl+KBPV+pNN4FUH+59yUIf1mIAiAI35mxarHQOBPowi/6hssMo8KIsbg4hwsXTmFhYQKFYgACEMcWjx6u448f/BlPnjzGnr1zOHnyGBbmp0AqV3M/M3+rkbz9H4+h7SAfpvfSloTnxgXulg3w7QMDXQYDg5FgYrKOs28s4/jxRUSRsxoYw0iAxV5C7y4uHjkFIHzZtyIIfymIAiAI3w3daOilXoI3B1YdSSwrCpgmpxpYXjmIlRNLiIoa0AQDwtZWF19evYkPP/wYgMGx5UNYOrwPYUFhGDTHvkyOXwX/ZPb7Fw3kezGeCUjM5faPbjaUBgZ+W3xAYAFYXJzD6dNHsHfvFMIAMLDUandLnV7v2Mzc/K+rMzNjkIBA4TVHFABB+E6MV4q1xhvM+mw/5oa1FmEELC3twYkThzE7OwalXJR7kjAePVrDlctf4f69+1hYmMbKyiGXGqhMVvSHfZncNMt/yPOW0TuPv7oe/2dtGTuUjJ0xf7m3lH4iu7abO6yUxfh4BceW9+ONN1dQqgQAGfTige4N4rlunLw7Ua2eGB8fr3xvb0wQ/gUiCoAgvDyqMsb7rQ3fsYyjiTEBFFCphDhx4hCWVw6gXNUuVQ1Au93Fjet38MXnV6GVxukzJ3Hw0F5UqwUQWVf5biSXPs/OHPud/BAKwPfrevjWV5caBnJ7B+yEyKtJTFBQft8Cg6gI7Ds4jZ+99wYmp+uIIoJlxnY3qa6ud46ON6d/Ozd3YBoyBwqvMTL4BeHlKRTDxnuDBKfimMYIjCgkLB6cx/ETS5ibH4dSfptby3h4/wk+v/QFHjx4hP37D+Ds2VOYmRmH1j4UjvJC3uZK4KbdDV0Eu/N9C38F+AqE3znTb9eAxK8PFlS5Z+lrAgMVq6waotsywYB1jMZ4CcdWDuLEyUOo1gsAGL1uoje3BhNBofo3RutlAFIiWHhtEQVAEF6OYq02uU9HxV9bxj5jjdJEGKuX8atfvoMjh/ehXAxA5Ez63XaMK5ev4qsvryGMApw7fwp7982hXI6g8rVuvHzbXYy/XtlrozaN5wcGprkS1u105KoDKoswBMYnSvjNX7+DhYUJhJECaQ2DoPB4rXXYGv7l0srKQcg8KLymyMAXhG+Pbjabs8VK6Tf92B5PElMnstRolLB8dBHnzqxgerIBTW4jnCRxG/5c/OxzrG2sY/HQXvz8/QsYn6hCabdfHtgOq9s9t3TfcyrjPfPcX4aiwPkqh/T8wECm3E+6VTEBSlsUy4STpw7h5OlDmJ5pgBQQx7FaXdsuRoXKz+u1qTONRqPxY74vQXhVkM0xBOHbUy4U6ksqKv3rfodnLRAWIoWFuTG8885p7Ns3g1IpBNjCWqDdHuDix1/g2le3EEURlk8cxuKhvSgWCSDrN8zJrWyfK/yfx1+GwP9Gnvc2s4DB9EGaUWGhA8LkdA3n3jqOGzcf4fGTbfQ7hvoJU7uXLJnEvjU9vXB5c3PzA7zK0ZPPJ++Z+aZP6EXb+yH5Np/xzkjX3f4K3wFRAL4/dn4JX/SL9E3RXcKrhZqampq1OjiPJDhnTFwmYmo0Sjh8ZA8uXDiNWqMMUgqWgV7f4uH9dXz80WVsrLdw5Ogiji8fQbkaQVGMnWl233bw/OVD+PZfCy8TfTGlIGScOLGEzy5ex/Xr93G/vwFmwuZWtx42i+frYxOXAVwGsP09X/wPwTA4w/2EcPO49n/9my/lz6dcYYmdbQ3/Fnc8z6N7TBdyj/s7GioOA1jQ+/rr5x0n7Bbt6sM/uxYo+2CYtsEwP9QASDCaQvLqp8C8gogC8N0huM+xUSw2apVKUAyCUhAEgUYIBMwEhMS5LxMRWUoSjkGcJIkxphu32+12t9vdBNDGdyr/JvzAFIOgfiLh8Je9gZk0xlBYUti7dwpvvHEMhw7vQRgBFgRrNTbWW/j04y9x7eoNVCtVnDh+DEtL+6H8/EXebw3gJyr48yqjQFDe9//NdQHcp6f9uUM3CcNgYX4C584t4/r1e1h9uoFel9Ht9pSpFQ8zhe/u37//97du3frkhTr66aBqtTo5NjYzowulSUJU6/T7laRnCn2OCzA2VKx8bYOAAEXGbxdlmZ1vyH0sNDSXWChAKRiCstjpfHKNqdxvR9G/NsU/xwBQeMZFZXO/FWyJWAGscq+3dii4LcjAwloiA0SGiAxgYk0cE3ESBKpfqhV7Wgd9WHQoaXXa7Y12t9vdbLfb23A6iMyhL4AoAN+NANXqWL1QOWh6djnUej8QjDF0ucc60oaImHQAKGLlvnzMzAY2QWSZjWEOBhalVqlSelAfK3xRKYZXrl///C7cIBZt9tVCVasT+y0Kb1kOTw2SPimtMTnRwPLyIZw4eRjFErmKfgD6vQR3bj/E7//bH9BqtfDm+XNYXj6GZqMGwOB58v5Fb/pPqS68yDV+9+t7ma2C00qKeauKQRBoHD1yAOfeWMFXV27g0YMWksRiY7NdAcfHJ2YWfrO+vn5za2trA6+m8Iias7PzsPp9o6ILxOERRjANohJrG2pbCAyBGKQAgKwmJgIxYMHk3Ex+kwnyRRUsvAuKYV20BSgrQgWvJgzvos3dUQYDbLPzrPsFgMDP2BkswK5lAKlWMbqrg0lvnAK5PZ6hiBisXbdkXaEMNgZaJYkJeyBqszVbhotPVDT2oKjqN+rj0fVKoXSn03n0+P79+5twlgKZR5+DKAAvjyqXy9NhVH23oMv/dhDQEc22QTFHsaVgoElpAiljEVgmxa6km9vPREGB2IKYoaylIAnCsF2ISneiYvhPBw8e/U/Xr39xEc9a2oSflnKp2rwwsLgQJzxuLVG5GOLQwb04dfIoFvZMZ0V/rNV4+nQDly9fwdWr1zE21sDxE0ewb/8cglCDlNmR4ucYnakUXiWrZn4jnp1X9H1bL9j/phdckA+vzYKIQcxgtmBF3opgMTlZw/Hlgzh14jB+v3UJ21sxuv2eKsVqjwprv2hOzv73QqHw8ZMnT1rf65v57uhSaXxaA/+zDct/2x7QQdtNGhaITMLaGCYvMYfDyZdGdn9BTMp9qOmYI2CoE5B3mKjR4UjuvjJyvgL/MdvsKPtTfZ4nhmODcg0x5awCPLyQbNwwj2gEBAVYcm/B9+USajQrQ6wG1pKCUUDCUP1AlbpRqLfDSD+y2nwFXf7w4MFjf0qSzt3bt29v4dW27PxkiALw8gSVqLKkVPBXyqpfVZiaESMgZuoahlWWigRMskXDWoTexmVBSKxGAoWEwD3F6BHQB6zpJHMmDOrzexYSa/t3b968+Riv5mrkdURF1eq+xOKCYTqaGITQCvV6EcvHFnH4yAHUaiWQMmALDAYxbt+6g08/uYROp4MLF87h8NFFjI1VnJKQbfYzJBVi7refMHdxgWdz5i4X+UNYBdhd3Eifz07yw3Pypo30PX2TgsD5RvGc9/ZCepAT/EPFySJVpIqFEAcPzOHtt0/j6tW76PVWMegn1Or1q+vrrWPNevM3BV24/+TJkw5ere9dKUa8v91V/1oX+VSScC1JjGImsqygdQgVKECRqyXhc0+z2EgG3LLb2QL8Ahvg3K6TxFm1RXckVRSctsBgX5RpxwigtHplGprgn/IVrBW7+hZpmSv4dgggJsrGipf0vk2nAJAlp8hh2CWDwJaRsAGM9a9RbBTDMGxi40Wl7JFQlY4XS6Xj8SD8v+t79vx56+7dV9Wy85MiCsDLE5IO9oWWTkeGpxo6xHRUIDIGT7tdPI1jTBUCnKqUsY8sSsZN+jErtGNGxwJ9IuoQYZUZN+NEb/a5plE6UioUt4DwPwFYh1gBXhWiRnXsrdjqUwnThCWmIGDsOzCL5ZVFzC2MQwduqrKWsPp0A1eufIFr165jbKyJM2eOY8+eaRQKqY96d4E4nF7dLLpT0P5UZv+vi1R1usyLWSmeqxBwrgna0ccOQ8noK2korHZeL40eVpoxNdXAqdNHsfzh51hbb+HpoI9eb6A3qTNVmW38lVW9PwB4glcrILDM4IXBwBzWMBUDpazV7q0phXKthmK5CB1ql1ZKnO2WmApW8p+TTUfWiMBnDP/kFQAvsr224AS3u1EWystum0luZh9+wJx99tov9q33OICHGzCkdRuGurA7j0BQRFCZwuGVEAbYEowxiOMBTBIjiRPYJKEkidFLEt2LTSUgLpcLwXS7Z/YVChHvKY1vd4Lgk5s3b35DfOLrhygAL8k4xnVgqR5aHq8lhvbXS1gZnwANYlxPHiPs93C0Ucbv5qZwrACUzAAAIWHCVmuAzUGCFhRaKsBNw0iersEwU0RU5QT7mM08gBsQBeBVICwWG3MqKP7GDNRBa02oFFCtRTh3fgVLR/eiVosAGIAJcQx8+eV1XPz0ErrdFt59922sLC9hrFEBqaHf9HmMhjS7yS+12tLIGT8urlcFSwQQg9hml/F8Af2iDJUd3qH4DN83QbGFyp51lQENmZFOM5mxo3UFi1IpxJ69U/j5+2/i+q272G610B8w9RJT2m71T0dK/2xp6fjtq1cvXX6pt/HDEChWBeggBENlApsI0AphMUKpWkapXERUDEAhIQxDaK2dosU8TIyknEHdurFIpLzAzqwGLjKA0rHqtINUWSBOrSoA0vgCIhArP0a8ksdpVYrUAkAjqQjs205HODP7OAMFlY6CzNxFgCWwAYwxGPQH6A8G6Hd76Lbb2N7aQrdjwAmBoahjbGSSzr65mfpvS6XC9Y2nT6/BzaWvhj/tFUEUgJeEXaiLUoAqgDEeasxEAWASbMJikxPMKcLhcoTFEkBxan0iJAlhC8A2A9uhBiHAZ2saj0wCaywNuoOC1mqsWq1Grdar5o587aBqtTpWKJV+0Y/1mcTYMbYWtXoJR5YW8MZbK5iZH0MQKoAYbAmb6218+tFl3L1zF/ML03jv5xcwPTOOIBquVlPL/tBnO9qpK2qT94vmzeo7JtHcGc9zC+y2an/RY8OO/aotXTD6FabmoXv5Gdi9l7ThvDl3pI/c8zYvzOFkQKo3cU787+xn+Fh503SuvCKlroEEpXKAs+eP4U8fHcST1XU8fLiBfn+gHj9JCvsXpn5Rq5QuAbgN4FX58rUjHTyMyuX7VhdKvZhLg4TBsARjsLG2jk6njWKl6H5KEYqlEgpRhCAIoLWG0gqKVFYrysn0VHsL3LFM3fRKGLkMPKdDsBfyDDWiYfkwTQIUE2xqvfEuCDXi1nlWTXTynUDQMDa/GZbbxpnIKQZsXdwBMYOsgtYBwoBhQ4N+EAA6LSftc0aYYRKLQAcLgQr2GBPUAaxBFIARRAF4SXx8rQXIKlhEBIScgOwABTtACQYVmyAyfUQJgKTnTJukoW0fVWucRktAVRNKbBGyxSCxZGysiVS5VCppUQB+csqFSnOxEFX+brur5tjaIAxBc7N1/Oy9s1g8NI9yLQI0w1qFuG9x5fMbuPbVLRAUllcOY+XEIRSrUa5IH4+YuzP3p/NnDidhGkrOVMBy+qKc/zaLuuZ0jTY8Rt4W/t2PuZk9W/d5kyx5e316/eSPIztvZxz/0Ibh+sj/n5qSsePsYZtZWzQUQIDCyAnpK8lmrgZmgMnCMiPQGtMzDZx/8zhu3nqA1dUWBomlhIm6fbNsLd5ZWlr68urVqx/h1RAYnXJZ36jVyv9PTOFvwgEtdnq22uuztgzY2FDf9BH3B+hstaAChSAKEYYhwjBCIQpRiEIEQQgdEFSgQJqgtQYUASoAlIImTkffcAmfWQFMFj/oMwmHumvO32/TkAFgOF4YmSvC3cucQ8sPccsEa60L3LQMYyysNWDLsNbCGIMkNjADi0E/hhk483+cDNCPB0jiGNY4JUUBCEhDa4bWuq9UEFNmehPyiALwkjCY4CyPVimFUAfZZEOwULAIFaBhnZ5gExekwwCsBVkLxS4XIDVravaZgkRKRzqyzmEs/HSoen1qDgjf6ifqzcRwFYpUfayMpSMLeOvtk2hOVEABYJkRDyyerm7jn/7pQ9y7+wCz81M4e/YUJqaaCEKXHpj6pjPYr4zYr7KcixXGT6b51CuVm1DTkQYMV9jPP+aOv/Ax3wzZdIVII3IVSM3JlFNKdloAchaL5/kEOPcaSi0KPlybssNQvg9N5JPcdmgIfqU40jDImbbT0ygVQgylGQVNWDm+hJUrN3HnzlPcu7uKxFhstLrNybHKm2OTc1dw9epVAFvPufofk1gp9UBr+j8sJ52J5tivS31eWd3sNbodVswAG4axDBP7DaRUH4o0tFbQihAoDZeWRO5voKDDAKQUoDVIK2hSzqmS/yzJ3STn9fEGehdfkC3oU6UsdTP4k4fjyvqx7e+LtfTMuLeWYYyB5VTgW3ASg63NnreWYRM45cBYsLGwSCtpun4UAVGouVIMk0JguiD6gmGuax1v49VQ5l4p4BzxygAAIABJREFURAF4OcjCKmjlHaIaOgzBugCjBkgogCUFaAVWCqwJMBrQBJgAljQSAANSSFQAqwIQaRAxlFJQSlMhiAqNKNKrX+9SlQH9w1IolZrHrNK/7AwwbZm1DhTm5qdw4uwRHDgyh6joUsyMVWht9/HV1Zu4ePESjLU4fOQwllcOI4qcSTpXCsr9ya2E2ACJAZI4Qb8fYxAbF16VswKk6dvgvG80PwSG6/OXGRqE4WpuqADkVAN61jwPuN34hiaM7OgOH0ee/Hne3kEMToPOdrwPDYIijWIxQhRp6JCg9Y7GmXMC//nvPVUECAbzc5M4c/oYrl+/h8ePV9HvWXT6fd2Li4f7A/3Ovn37Prh9+/Y/P/8T+/F49OhR59GjR59OT88Hs9ML46VaMG1VWOt3t5XJl0BmcnF51sKShY0tYjY+5S9V6ABogLQP5CPlFANfqiSvSGZaGilnfod3BVD+89/h09rpn7LuV/ovW5WzCHjrDAPWOgWAmZy7xrL7odyYSv0XNnePVfpdMChEEU9O1pPZifpmu7X2uUkGf9/v9D5uNBrb9+7dk/lyB6IAjJJauHbuO5of0gxA9YtolpVuWOhibBS6UNiyLsWvhRA9BGhBYRuELitoctU6GRpdJNgAYRsaLYqwCY2eCpAQw0IRkQ4bjbHphHi+XJ5MmJlKJfct73aJibq2o5RBqxXDFQzqQ1Jcvm+o2GjMGq3fYNLnY2sCUoRKpYDFpb04efoYKrUIFFgwE5LY4tGjNXzwwUd4+vQplpYO4vipZUxNTwwd2OTCoIZmc+0mPsPodPpYW9vCk0drWN/YQqfTQ2Ksk/Uqe3mWFmX9wWxSBkBZfDXnfvKefXrmWH5GzPz63k1BdvQ5EHkFIDf5s1MAhq2lL9K5br1XOTM3sF+1EZy/Hk74pxN95oNwbSoiRDpCo1nDxFQT45MNjE1UobVzhaS9U6pLQIF3SftOo+IJFuAElXIBR4/uw8nTh3D50hd4+rgHaxnbrX5TA6emp/e+f/v27ct4NYpyRc1mc6ZQqU10+p3IqgoHOsr5hSizv2dCMlXK0hV5fhozFmzS+5AAcBsvuXbsDsUSw9dms6L1AyYNKIAfFjklgzE0RaXnI6dhZn0oP8j9mKV0U6vAn8NDxYK8ikK5VE/2789aVMpFzM1OxYsL4w+uX3/69w/vPfrPd+5cvwogfsnP/S8aUQAcYb1er4WVsZlAR3VKdImVCYBR66izUioTJyAT9/fHrE8RU33LArfaPfRigun18TgG1jnAjb7FJxtddCJGycQg1hiwwmonxkbfogNGe6BwnyzuxcCm1TB9BjpJqTZRu0CqbxsT40/YQilibQEulMhY5qTMtqfr0y0d6MdRke5iMHh48+bNLYgi8H1RLESN87GxF2KmaUtAMSIcXJzHmbPHcODgPCjNgYbC5sY2vrhyDR/84U8gYhw/eRSHDy8iKgRwRu3hbeE0iIqBJAHWV9u4evU2PvrzZ7h+9SZW1zbQ7nSRmATMfoGTyk6/BLe5+TiVyWlA1ejSS+X+p2eOORnhV3jOsZVZHcikDaetElgNr99Z32kk0Gu0r/wVWmirvSUkTUdzCoCrUeOizr1FH2mn7tUKYVDAWLOOvQfmcGxlCW+cP4m5uXHoEBhNJct1/QxDywOTAakYM3MNnDixhIvHD+KDrSvotBm9/kAl5eLeqDz2m4WFhX9IkuTqo0eP2s9r9UegWK/X9+qo+m90UPr147XusV6/P9mLSRtLXgDuWLNwTmvkHR9MZq0xQ6Gt4JUGGhXGI+SVgPSxzt9ijPiBMn3Dp70yDc/lfDteiVD+ibSmQH6bR+UVxJENn3LH2ADKbfecxMY8fPK4v7nR7g54oJrNZrixsZH/YggeUQCAsFhsziOqvauD4vuKCnOqENRIKQ1OXVh+3UNgMNtAWwsV1vqDZK4X23LfAv2tNu6gCzYW/ZgxQAGmzRg8WMM0xSiwAbMrANRJCF2j0IdCV/WwgRAPEmBTaZhOQptPt4uVQXLKJthLUX0A45aNPiiLlWWrAKM194NArStlLuow+sdDhw59cO3atSeQgf5dUfX61IJWxXdi1itxokLSFrV6AadOL+H48YOo1UtQygXzJX2Le3ce4+Inn+PxoydYWV7C8vIhTM+MQamhj9JNXW41xKxhmbC21sLHH32J//KPf8SnH1/G9nYHxrhqgqSRM/f7Aiojq+MUQlaWdYRU2PvV9ogC4I5xKnFJw21JnA4eC2LlTb5eaI6sCtPl9mgcwPBZGio6vl/FGpQWpk0XgKz9yt2vEp8pJkSwVsEmhDv6Ca5ff4ibNx5ia7ODX/32HUxNN6Ajn4Hhu3uu/M9WmF6tZ4NCQePA/hm8+eZJXPviHpLBNuIBU6vdrz5+un5sambhd9v99v/+6NGj6/iJlOvx8fEpCkrvkC7/h82tZLGX6OogQWCtJnBIo1tE7xTctONnx86THhVo6CAYulFSu3z+3KwoEDD8KHIWAJuu1LOUjZyykd7XXHtpZgG0VwDggv4S42IZ0vZT5WGYSDV8L8zIlAGlsdFqYXC7VyxHvFgOw39Xq05OVAuV/2ujUPgYP60S90ryuisAqlKpTASF+lsqKP4vg1ifANBQikMiq9JUluwrQwCD2ViGNaQSo5Uh6IFS6BoLzdYNxSAAWMMoi9gY3CFCAOWCuwgwpBFrjb4FOolFlxgdFWCgFVkLpk6su2ybmlB3IbND8x2x+5LAe8q0TvqFEPvLhbBZLEUE4B/gNhQSXp5CWCy9k5B6IzZqmplVFBD27pvCiZOHsGfvNIJAAWzcrnJrW7j65TVc/eoaKqUy3n77HA4e2oNSOQRotOZ/3vDe7zOuXLmJ/++//gl//KeLePJkDYWogLHxBhrNGorFEERpHD38YpyyZCdX3MWrFdb4x/lkq7y5n0aOpW0O4xIUrHUWBzdnO0WBMjNr2mfaghcGlC7C0qyE4W+bsxS479JwZZkqAMR+8velYvK+YZcCRogN0NpsY2trG0+ebKLT7WEQD1CplfCz985iZroJUpRZZL5OBRgVfhZaKUxNNXD61DF8cvQLdFpfYW2th143DjaDwdTEWPNv44Q/bTabTzc2Nja+puEfjEKhOh1ExTMDUzrS7tpKPwFZdrFHSPf++XrNJxPeQytATtHShEKphGq1Cq2dSCBfTZG968ZVEEwjBIZjkr0SmI/yd0HQeUGPrKYA5U01DGdt8EWLUu9Du9VGe6uzo17Wzg2G0mM88nw8SGg7HgQDjSaX9alGIyrpUD8dX39yew3oQiykI7zuCkBUro8fMSj+JjHRz/oJV0hDayJoKDC7NCKblqNk+MHuJ76IoYIAIAWDNC3KfQU0AboUQJU1WMNHq8KZWk0Am1j0uwNsdfpIKIRV2lfvYgIxYmYkbDT8RJ9+SdJ8XLYAGwPbj3UpUge01lpp1VlYOHDn3r2bnyF17AnflrBYbMyqoPSvTExL1pqi1kCtUsKZM0extLQX9XoZSFNABsCdW3dx+dJlrK+tY2npEN44dxrT02NQo7bxDAbAhrG10cEnf76Ejz+6hMeP10DQOHBgHw4c3Iup2XGUys7Hy1k0vhPJNByMyFZk1sUigHhEDlBurh2xEGM0PY+hwJz4RV/6TM4UzENL7DDtMH8srU/j3ATKuqIzWUnaHR8Fw2URaKNhlVv9UxrNn7M0WBBiw2itbePu/Ye4ffseNjbWceXzayAaYP++WTQbVRSLGvrrBOAzN8GdrIhRKRWweGAev/j5m7h35zG2N/uIY1C3a4rbrfiEpuDdmZk9tzY2NjaffSc/POVyWEisrnOMkC3nLCu7sYulOzvVvy61KmU338WlaEXQaRlh8oGrIJ/fn6p/fsz519q09HDuOcV51TTtYqigEFILDCEtB5zZe4igVKoU7vJRP2P5St9y6vJQsNZQwkZ1u0mpXouWSNEic9gAcP85H9pry+usAKhSaWKCUTgHDt7rJ6gZVqiUq6jUKghCDWst0rraz5o/Hb4ch5+Y2bvTCIVQY/+eGSzOT6FeKeY0YoXEAKsbLdx9+Bj27kMYFYJJwZJyxS6IYdnlxKa7c5HyXyC/aYZNDAbdHlpb29SL4yDsmYUw0O9Mzkxfb7XWb21ubsoGGN8eqtVq9UK5ciGx6pyxPMFsqFSMsG/fNC5cOI25hUkEgXc7MqG93cWlS5/j6tVrKJeLuHDhDczvmUWhGOJ55lYwkCQWjx+u4epXN/HowVMEOsLk5CTOv3kaBw4uoNasQIXudOsVADeHksvVZmQKodNLybkHnJUq61dlefa5/H4gS55Kr244Bac1CnJWp1x7xCoLEnzmWFrnTQHOlJW6JtgrByqd9/2rCWQJlkymOBMNYwqckuBWhckgxvz9WQShxpXP+1hfX8UHf/gQv/vdr3Hw4B4Ui9WvXwHvvNE5k3moGOONMt599yz++cNP8fRJC0+f9hEPYv3k8Vptfrb5frXRvAhXmfNHLxEcx/GmBd3WFHQDzWFsmQzbodsk89m/qOUjPc+7giyj3+liMx74FMChwgliqNQCkAUZIhO4lqwvIkRwsdM8EpgK+Cl0x8ZXbipLx2TOesGEODa+SmHeapV3Y+3y1nJvnwC3IZQCtFZxoFWs3C5dwg5eZwUgiiK9Esd03oD2GiYUq1VMz8+hOdlAEGlYtsNiKFk0Ko2ujdJdt/yuWsoyNAH1chEXzp/FhbOnMDfZdJq1p5cY3LjzAH/65DPEH34EowK4EqvDCFe2wyna1cb2j7xvzhiLdquDh/cforW6gW7fBKUi7ddB+V9NTU39QSl1eX19ffMn+Fz/JVNQhcIBraO/6w7svDEmDEOFyck63rpwCkuH9qBa8SV/LcMYwu2bd3Hl0ldot9o4vryM82+dQa1WgsoV/UHuj4NgEuDxo3Wsr2+j149Rrzdw4tRxHDy0iHqjCBU5symzW5m5lzHSaG7FKnNPwU+i6V5uTth7Eeu3gSdYt1oDcpXcKNvuNRO6uetMW/Nqrj82zDTISr7mKu4xyE34ijI3QTp5a9a+z7yKwlAcZB06j7Ar7MPKCRLNjDCKsHf/HDY3WthY38LTp4+RmASPn2yg0+1hnKrZ9Yx84CNyj5DLVs+9D4Mw0Jida+LC26fw4P4GWts30esm6PQsYoNjzPzm4uLiZzdu3PgUPzK3b99+MDe394/VauNTFekTaJlGp2+1dW4aGq19nBPeIzeTck8ThtH5Ln7CWIvBwJdUptT2nisbDDhLwcg44UznAwhk3YZDwNBBADj9hL0y4Ssy+TaGkns4O7qize6cFyyDwsMHREAhDLhWLppKEb1avXKlGKkvWtvl1dVVMf/v5HVVAFSpND6pC9V3Y4SnB0aXdRTR+PQUahMNFOtFF4CFVAkmv4hhl/YPdhNmGs3sv3/kzbMBM0rVIqZmxrFv3zzmpyYQeGFgCegnBgNYXL9/B2E1dCYvX/3adeonQMAJfD/FWkJmZWAwgkIAYxMkvT71Wi212e7WmOPlsfr4X09E0db6+nob4gp4UVSx2JxRHF0YGHrHJqamialZL+LQ4izeffcMJsar0AEAZlhj0d7q4+OPLuLunQcYG2vi9BvHsXffHAqF/IpMDavdpStrX/Vsu9VGrz9AYi2iUog9++dRrpShA5fGZi0wGCSIB9a7ftivtoZzae7ysdvqaLieGxYhSoP28gunoZWYsldp34GlVBklaJ/znwafA4D2D+zoy72yklMU/GYxRDY7lplus+tlp9yQhY40gkhDa6dUFEsRZmanMDU1CWMMjFHY3Oyg2xt4FcVkNovRvYa80B+JIM/DgGKEBcbps0fx5Re3ce/eYzx8sEHGAE9Xt2rNZunc+NT8pRs3blzDjx9js7Wx0flM643/bf7A0f8VD1vHB6vd2sAwDYPggBGL0ws7KpzFJigEKBTC7J65e+jclspPhiqtPunnHzBnpX/d4seNe0vpXfcKp07r/DurZrZtsF/MpEkIIIJlIIkNkjgfz7Hbqn+nRYMBtogCjYmJqt03O94ltC7Fcec/rj5Z+8O1a9d+EvfNq87rqgCUw1LhhOXwnGXaS0qrcr2GsalxlGoFUEAj81K6lkl9rE6DTlc/ueFJlH0HSROiKECxEKFYCKF9MBcTAwEhKgTQkQIH7lg+aCZVzhWGXzgAUGSz7yaRQkgh6mN1tDZbiAcxer1OECrMNJv1Xynuf16r1R5tb28//WE/yr8Uxqu1Zm0FiH7dSzALcBAGRPPz4zh9dglHluZRLBKU94v2OgPcunEXn3z0Gfq9PpaPHcbxlSMoVyMolWSrotHJK91QxSl4SZIgsU6JVAGhXC1DBc4cag3QavVw7/5jbKy3YBK/lavySqGfp58dhaOT5XAdly7+ciuwHee5p4cSXPmglnQyJ4wKe7vTegBn6nVfE8qsEJxVhfO1C3KrRGKdZYfBK0jEBKUZYxM1TE+PYXyiAeWzzUqFCKViwe8Mp9HvJUji1Lr7dfN7fuXv1YSswiG7VS8BcwuTOHXmKK7fuIfVtXX0O0CnO9CVauFwbMK3Fw4c+PDezZuffENn3zdJt7u6vb7NN+eALZDXdHZewTPHeMcTu7kI3D0KwgDlasVVCQQyDdOrsACp4XyUNU0+zsPbElLBjtRSNezSKWhp7YBcvQrOtgd28VaGsb3dxnbc3t2CsSvD84JAo1ot2/GJZmt9dfPi9tbWn69cunQXUgdgV15HBUAXx8bGw0L03iBRRxJWlaAUoTnZRLlehg41WA0NlKlZc+hDzTma/J8sJ5u9MYtcEI1Kq6Glc25WkMNvzEnWKxrpBJnNgcMuCH4i9e4AyoXXaEKhXEBzYgy9Toc2Bz30DUqt9uBYMYjent+/dO2Lzz5ah8QCfBPh1FTxkOXoXWvDt5LEREQu7e/Q4T04e+YYxsYiaL9AMoaxtraNf/7zx7hx/RZmpqZxfOUY9u6bg1Jm93kWXuDsMg9nqc5K+Rx5Qq87wL07j/HhhxexutZCkphMwAJuQ5RhejflpncaadfVZ/cBqEwApSuwvLTIG2CHc7drerhBS17NGHp5054zM5jL57fKKwPPysnUR+wuR/sIcRqmOIKhNDA93cDSkb04XVlGqRJmBmHK1Q9mi5EMyGEZ23y/Xy+r3efqLASFcojDKwdw8uZhfHn1Bh71W0ispXYnHleBPj05MfvzezdvfglXHOjHMinrUmm8UQgrpx8+XJ1ptUzBJHbov6FdBGVqMRo+Mfwzcsvc3GJMjEG/B63VMBCT2G/+415IpDMVwAV+poqks4KqnCUiX+4/PcddXn7+9OOAvWqsFKyBKxuQ3WKLzBXwXCXAZu8nMRbb2x168Hg1MN3BWByb5sTERHF1dfXrNIjXltdNASAAFa2iw6DobcOYhVKqVCmhOdFAEKlcQEtuIs1eunOqTJc+6RmuBpliBc1puFZutUXw22IOV0qjbe5cM3L2l0euwm+7SQCFGtVmFbXtOtrtFvqdnlrfbtfmJqpvFcPwUwBXAfwk6Uv/QqBSqTQdFCrv9wfh+/0BzSQWKBYJexamceL4QSwd2oMgtCByQrfT6eP2rfv44I//jH6/h6XDizi2vIRavQKVrXyenW9GAknTG52aXFPhCbcxSmu7h9s3HuDip1fR6xkwKSitvHXAwiTsqqGmK3byj3cIXDdKbU559XUAspq/GBmAz8rr58m4vKDN1xpwY9vFHuTLHz/bR5ZCCB7uCucvkRTj8ZM1xNbiwMEDKJbDZyz3SqX57+4n24sj+0zTS8oFlD1XF/BVDrXFzMIYVk4dwsef7sHT1S8R9yy2O72AAtpfqlR/NT09/V8fP378Y7oCigD2GEP/4+ra1qF+EpaMUW4lPbI3Qv5G7lSE8s/545myYBH3utgc9JCmmQ7N/Na7ITFUANKFTtZD5gTwR2y2YMruSbazsLMmuDHrBHda+ImUgmUFkxhfU2C4YHquVp2usPxGAP1+jIeP1/X29lZzbrzy82JU3ZydXXhSKBTW79+/33mhT/s14nVTAHStVpvVTD8bxFg0VpWjagn18SbK1bL3+/NzxlvuAA+PjaxwUk0W8EVURl+drtytn/1dzEAudGk3k17aT3ZKqlRw9nxUCNAYa6DT7mG1+wjJAEF/YA8S89n9+5c+vnXr6se7tC4AQbVaHS+WJ37JKP01K5yIEWvSjOZYGSdPLmFleQnNsTJ8fgaMAR4/WsWlS1dw6+YdzM5MYXnlMGbnJ4cp2QCGa56dPH8ys2BXDY2ATm+AjY022u0+CBHK1RpK1QqUBrq9PrY22rCxdbsGAb7NYRBWdghwE27Wpb/I1OwAjJybt0C9OPllZVod8dm2M30598psXOcCHF0mrMX29gBr6y202gPM5FMS4QXQiHYxdFO8zFAfugMsikWNfftncPbcCq5cuo0N20MSG7S6gwZWt09Mzu7/H4Jy8/+8f/PLa/hxTMvRwCZjSS/eqyIuppmVzyqZO1b8I/EVuZswouUpgNx2wUGg/dzFOwYC+8xBlcVD7U7ah8rmxbSSBOnhOcNYJyfg2SuySmuQTV1L/odz7e5iTXrGZAUFay16fROsbrTHF6Yr56vlwkerq52LcHUAZB7M8TopAAQ0q0GhcphV4f0kwbgKA11r1NEYG4MKAlj2W14+U9qMRr9sDHAaEJNbsmdWN3b/ZFtZ+h2tmH1ak2FntrTIAm7zSoBKhQcBw53YUv+aVwdy/SqlUa5W0BxrUnuzhUGrrTa3ug3VLJ6empl/a3Pz6Y2fKof5FYQAhM1ms1wqNeYSFbylqPwfOgN7pp+YGmtDxbLCyokDOH/hOA4cmkNYIFi/yG23e7h29SY+/egSkr7ByRPHcXBpP6q1Egg+bTQT/n5lku8Zz5lAMwHsFA1rGUliwQYgpdAcm8DEzCQoVNhut9Ht34VJOn6cpCZ9jWF0dw7erbb7zu0udjEXvzDpYMwrN7spzF9HzqzPGkACNjFM4jJewEO7XBpsm+6rQMT+i2T865FZFEZ6yFayo8eHwt9dhtaM6ekGzpxdxj9/cAmXL9/G+lqPBnEcDPp6Jhwf+5/KJbsxN7efHjy4dRs/fIEZGwRBUiwVB7pQtp0eozdA7uPeYXXaOXc9o4HtuCEqQFSIUK2WoCm1xuTmwNR1xcPP/pk20/+yAkNuKLraj7nTQVk5a6hcQSHr7qVloLXdRifpDBtJX5++31Ez6fAy2CmJREwEZqVI61AXoVQxDPthrhXB8yooAH7XB+ipqSnNzGStpWaz6Yx3Nr//WNP/3YB6XpUVj7V1AgClthgAOh0VxXHvYEzhO8aGKwmjXCqUqFSuIgwKSAaJjyK2OR9jijN9DY9SNiFlfk52BTCUX4n09ADbrQ6erm24L5XXvC0BA8PYWNtGZ7uHpJcgSau9+cHulGU73NsjW9uo4VVQmhUAkFUgVigWSqhUauhttak3sGGc0KHYqvfm5vZeW1w8flmp3qDXi6xS2jeye5ag1jp7qyO+g+/oSGj622eM+bYS5gVoZI+sNWQqo33UAcRxQbXbW9GTzdVxrYsHdFQ8x6zf7/b5RD+Om5ZMUK4F2LtvEu/+/CyOrRxwq38FABpxAty9+xAXP/0c9+7cx8z0DM6eO4X5+SmEoS9Hm/XIGNmwBBia64dn7DIduXHitsYd7n5WKpdQadSBkMChho5Cv5c7oIIQSqcr+1x/2YyZ00yzIIRcidXUTE47rnFEiO4wxWbnYsf5Q9IMlrx1YeQUHqpKaXwEW8AM0r7UUPDnrAd5d9gOEQ/ONlDePSvi68hUbLKolEMcWJzFe794E5vbHXS6D9DtGOr0BqXHq9vL5WLx35bq4/VZpj+Uy+UbUVRt93oDo9QWK6V4LdfueO5xfj6z1pK1NWo0ds5zgFKKNzcBpbZ5ezupVOo1bjQnV1WhPnv/4VY0WG+RtX6M5VMv/Gp65NPOBlp+XPjP15f+tez870QMaD/LZJlIrk3yC5vh5/tsnYusIqAv/JOJeIKrFsns61gMC1ylQ5bTjAZWub9pw7mxtOvMP7QWKK1RKhUwPz9lq1Vqs+1QoVAbW1paiguFgnGzwYuwBaUUb2vN2HAyRynFGxsbHEWRuX//voHLsvoXG2P1UykA6QwUAZV6FNF4tVoeC8NCFToohopCS4UgVEppDWLFpL1YJAs2qIHIWsByTMQw3g6qNYWsiJVSWnsBMCixJcvlRlTqdIvLg575+SDGpGGlwIRBb4CNpxtg5aKsXdDTaC1rQhr8kjcwDge4+4+cIAZDw6BXivDZp1eQdHto1kogpIF/gGHC49V1fPnVNaw+XIOl0BXP9PP0cCJKu8yrvsPveLa3hiWQBeJBAliCZUJsrGr1BpNRFL41NT5ngij4dNAL2wWVDGASJgIbU/QGCDe9GgCwBtZadp8zUAJg/d6bupzdPjYvNOQ5SxvXAOI4/UanNdv0C6T65k8Y7VQrDYYbG0pZYk77U8SpdISFYibLpMKiDkuqUakOaKbTjw90+3TUkjrY6/dChlXlisa+/RN4//1zePOtE5iZG0cQ+Fr3Fuhs93Hpkyu4fPELAApvvHEGh48cQr1RAWWBozsnWSA/a2XiNIvk3205M5w401KrKlBQIcGGBAoVoJ1iEBQClGpVlKoVb7nasemQr7KW+cUtu6p9qSrphxmUq3mhSMFCg9P6MpkVKm3bKTrZ92Goj3p9YfhestDENOsgW13m3me6Kme3JfKgH2P1wTr+f/be7E+O40gT/Mw9jjwq6y7cJwneh0BRFFtqqY/p3d/2/mZmdx/3bf/EfZuH7m31zPT0drdalMRDEm8SBAEQQKHuIzMj3G0e3M3dIzILKIAAWCRgZKEqIyM8PDzczT4zt8PlvKAgfNy56fikjRAaQvAByNlPEgCnCQuLM/j5z9/AtWvXsbuzj6tfrWI0HKs7a5t9Mzf4qQbm887cC73ezKddInScAAAgAElEQVR5bm9C0x7X3aqyxg4k6QLXbqdbA1wzATlBg5RSKmf3j7VKsSqVVm5dGAJba7k7Y2qu+2ZhKcsHg/6pleMnFWU9u7U95o3NPbIsAMAl4JkU/unvdD62xs4w6mGFHVO7jRZNkH38MOicFn3y1ibYg9uV08ISUJ5fUdJHIPhnhK0Fjbqq0ShmJI2JCZXQnAyS1dADFE0Kg8EcTp48yYr2y72t6sX+7KyFqTehAAWLmFzjADKWre1xzdb26tpU/VnDdW1sZet+f3Y0Go13+gsL6zzSq/0+bd2+fXsIx6C+VxaG7wIAEIDu3Nzc8X5/8dL+mC9aY85bheOVzeeJqWcVSmVNXhFrlwGXCKgFfbJlw8QOABiXLtwN+phpRFCkFRGTUmCwZWuYLSnTqYw6ZiwfN8ZmDGC4N0Rd3wbdWUNUM2wMW/LzX0E8lN1EDVhdxcVBcFq403oM8oyxubqKP7z3LspCw+WN904vpLA3rLC2tY07d7bAnMGS9kwPLg83iVOT61MKAoIHttfQlEfPbNmFizFQW6at3WGutLrQ65THsD/6ZT0e7dWmqsCWwRaWIRmOHCAnuD6CXX4jkRGWWZF/WB/rC+aGzZM9hHCFPRqC2okQAhSBmJi8JYNUkrx1mv20KTLBIniiXlC59EuUkc/DRCDvtx7vAwITESulTF7X3BtbmqkqdKvKZIZqAhv0BhoXLi7jz3/5Ov7Tf/wlLpw7hm43c+6WFrA14Ztrq3jvdx/imxu3ceGZ8/jFX/wcKysLyHMFUn7tpw5obpIkw9B6uPAS6QC2IaGjLuWq7JNLNT0ooOgWWFiZx9LxFVecKAEgqee+JmfZYrZglcNISllySaaUMq7gGhQsa9SWAgCQ+R6qAPr3EM3BYp9qx9dTOObyv1gHlBq5hAXjKtiasb2xh7Wbd6YI+9Ta0DTZuzHWbu7BCa9p1Db9p62mB9gj67LUuHDxGP76r97CeH+Mavgern69RqYmbGxuD4os+1G/k72wN6429djcGddmhy2PjTNi+nWlSCkANZO1TESGqIYCWaVAiiqllYImqomIFMjNOGZwbUzFBrXWtcLeuJNtbJ8kPSqGwyGYDYIXpfJOcyx6VdtqcxCJosOwlcG49sJY+I4oQxPDKQAAmCrz2oMa3lFrfhC56xu5DLLA6ijhe8FvwOehaPBEQbL+3RMTTGWwsbmt2Oyd3t/Z/Zu9Yf0226oCExHVYRepHQ8T+8xsma211lhYY6w11toalipj9J7hfKvM57+ZWexe6XeLz3vzxz+/8sm168D61rTmjio9bgCgBoPBIuWzl/Ks+HPLxf+itX7OcrVgmcuxIcVsHcthkMw8WbjMTrCQeKaS8/y0SpKVshi2xMHUHSUwW6aalaotlNNyLOrxCPV45Oc8+XAkL/W9cEVDU5M4ZkrC+hDTsbHkQ69Bqsbe7jpuXFdOiLBpiHILoLKuHKxbTJ55Wa9pJQCAJZ2qv3tYYUGqwml2AEgpF6tODLYWm9s72XB3d5ApNQM2ASt5EQLFDCny4TK0WYjbb5KhO4kPV4il3JKZLu8jMIQW16CAJ/z3vvxXwi3SJ5QWVGAAiNps4yrHjBp6DsWrIyNjEGuyxsJYJmYmJkKWMZYWZnD24greevtl/O3f/gyXLh1Hrl1xGfba5XBY44P3PsZXX15Dv9fDK6+9hBdeeBadbu6EWoPppU9yCGJCOyFOaEdFj2qRmyypqZmhNKHsZhgMOs6wEpLsOJaZgzA7N4N+V0OT80cZWoW19S2MRiOUZYG52Rn0usppRlZjOGSsb+6gsuw3xRBCvlJx7H4kOyUCEE4pjYIhAKxM1OzhQrwkDtzWjPGodj6LlpMWyK+F5ptnrzE6wZ/ed9pYNka11cfpZxAxOiXhjcvPgccGtqpR1b/H1kaF0X6F2hi9s1/1dvdH3Uyp41ZZ67YAXXii6NGufQsrRXLaSWwYxGFjnRjaPbMxjhGRUtD7hu5s7lNdGTWqCNa6sDxQ1uRXacRDAgAOmonhvSBpIwx1ygtbfW6s0tZ36fAH4Zz+pnhPSEpjoTqMl3DbEIbdeP/+2RrSW4EIMPUYd1a/wdb2TaWUGRCbGZBlma+Wnck05B+AvBLP0yi5AyXLDgBYgZkYrG2hs4pUuW04+7jI6J8vXjr+P7ar2fdXr1xZxfck78DjBACq3+8fU/nMn2dF/z9Yzn++O8IZw+iz1TkpJjfv/SshyXwepzCHr8nPUycAlaJYcd3PWaVdeZNQ1UoTFIh0Isgd0ndKMIEBJe53HCalFMOg1Mzoc283pnPQ5jwSJw2lGErJOvL39LNNEaHICHkuwYPiaOOZKKVCV4QaRGmCpB4OwtlrA84PRnl07RIIK3gGI3LXC3JZ1wTH4BXJQvMZ1Si2r8IyoMQqL8BMxkxQ/qTmERZ8Y4/av4sWdwrvnASgSF/ctNBAyGYXtYu0AYZPQO67LNcqlMjA1kBpoNvNMb84g9dffw6X33wRL718HufPLyPPaxArKFZg1tgf1/j62m387nfvYXNzC5eefxaXL7+GwWwHStnIJMNz3F0ABWqY/xMJP5Xc27bsc60H66sDjKRc7n1LjqG6rSSLTqnxxo+ewfkzyyhyRmUMbtwZ4l9+/Vt88806+jM9XP7Rczh3Zh55xjBG4+b1Tfzmd3/A6sa+53rK7ax7jpnCKzfcDhC6eZAAP5lyiG+cyfq9YHl5NhrSFIO08SPo3qErkOXvkw7PhDYf1/XhFLAmoEmPivFL+9v0exleeeUiQMDsbB/vvfsJbn6zht2dMdU1yIJc8SMGs7xDJatT+yx3GiALZYGo2MTxMYh5RmS8yIckkxfGFjU4c0xbnlSlwpMF+FFTaDfgPDceP8L4kLfPO1X6z+l6bSN0Px9CF/yzpWkmuPFE7PmNAPP0vn4zUs4JCYKixbMdcdV+FllPSpCMMoCyDhVAO+AshYfc4JPMQ4nZSh0Wk5QFnnUxjPG1OSxgrSnN1qij87rX7RUne5255+ay8h87Z7Jfff31Z18DGKE9wY4YPS4AQMDCQOXdP7NU/l/jGj+zzGcqg5yIkBc5FaVGWWrojEANhyQhpwsqBehMIc8USCkQKVilMSbCkBSYGZqBgi0KMpSxhYYzi1svvGOwEAX4pxheePrJL+jX39sJQvgMZxQFMTgKxzATJR2g24lmz6hd9jQ/7xWJkA5PKJECMvGUjY6GNgEA0vcwQdl7fyvf97APnCw8AGSNn82J4OH4JykR6DYBAHIPAQPuIgeMRHh7/4Z4csIsyJuWBVw0zkzGDDFm2MtTQ74QiYxb4GtNS4AlQFkdTOXxmQPsABGgdYZunqEsFAazXZw6uYxz50/gxZeexfkLxzC/2EOnCygSsyShrizu3NnGO++8j08+/QyzswO89vpLuPTceeQFxb31hhZ2ME3nBjR5UmuI5AzF8YcmTuYgVNw2TI0sVzh9agHPP3cSnZJRW0Z5dQu/f5dg7RBlAZw9vYQXnzuOogBMrdDNMnz0UYa1LQOqtR/3ZH+8MXWEy7sOWT/lFEfWnr4N4bqxdLGNtpqQOChl9C70jDkCzeRpW2OaAObw7UF0MF9urmYLpYHFpR5+9PolLC7M4rlL5/H5F9dw7eptrK5tYXd/hGpkUNWVc2P3vEazt1+F3BBOqFmyEPjO5MBcTTbwswkv/RAiCcCqsOdJ0NA+QFVOAxCAfPNRE3A04eQct5qIVQAc4gQoTYRl7c9ztRoQwVwre6+Dd/5QMi9CX8j5RMk2q7tRfBbx/xD9ptHrFIyEY5IPwt3ZOkto2Plh5rit6p/P8W4bQIklgVCUtu1LsFiMhjVGwwrjkcF4XNO4qgo2Jq/BMwzMD7q9lTzXxTPFi3/3+ecfXoEDAUeWHhcA6PTms2fysvsfh5X+panVactWk1bozXSwvDKPpeVZzM52UeQKsa53YN8AnDaQ5xr9mS4G/Z5XODUqlWE701g1jKqqUTJjoAmzOaMHi9zUPmzPSRHWXiDZqP07BoSALG0AAIyQaISFbflEKh4lq6kzMzIyMS8FQcZO2IozVpzZHNa+LCzBQVIlkKc6jcUJ687hyXMYIGt9n10bEV+1N/maq8vJNW+QY8f0HdNOynay8XvF0mm/sJV35oKPc4dklZ+8I3kTniQesWCQFfQP740fRiewe4YrKMMURtm3Ge+iNCHLNPpliX6vwPz8AMdPLGHl+CIWFmbQ6SiXxQ9jSA50toytrV189ulX+B//9K/Y3tnG23/2Fl59/UUsLg5Ayghn8Nzq7iJHBtAx29R06sZFtJ4pF/n/BSC5RFPR+pq8pwAgnUOrUjU6JaHX0yg7DGuBTqmQqRqwFTRZdLs5+l2NTgFYo9HvaBTKQjOjZtHGAZv0Ld2OCHOd0rwY8eTm+47ALLwj33YQ77L0RPtre7WHlqbnWojuKwe9j/ZVrfNESwzPZqAzjfmFHvoz53Hq9DG8ensDN26s4vbtdWxsbWNvd4y6rsA+xNfh8WjETkkAAOAAgGKGIZfYKGSLDP0UpCf79TF8k5CE2SHKdcnkdzAEmgIAPBtSHBULMMf3TOlbg1eEIp+aBqiE34VhRQsAwPoyw3A1JqQvaZscnVZdlxKQm1zh1EYBADJyfutv2jOH7V4FkPVgTf6LSaXCPRiw1mB/f4ytjV2s3dnCjRt3cGd1AzvDivb2h7m1fEyT7s/1Ozm6dvvUqVP7169fv44jHCXwOACAXlxcXKa8+wtL+S+Y6YQFtM415hf6uHDhJC4+dw4nT69gfraLIgPCy0reAbMr7zgz28exlUUsLywAZGF1hj2d4ToTPt4bYmd/D7MEnOkVONUrsMAGBTuNTgCAbC4we7Qte+ze7M7CSSHatKTHhF8JPjxJBE5rwUa2JFnXBMZwABlEylkBoEI4jF+3kWw050WB4a6ZJGkjnbiJLuNmcNIHFdMQN7B6ei3HViiGmZEX5YQMIVuX9QAgAW/wWywKsWytyCsFNJckO40mCC+23qLo/RRVCgCECXJkfz6nvDvm48GhI6AiQGtCkSkUZYaiyJDnGbLcC1YfKy/WGQuFUWVx9etv8M5v3sWfPvwQx4+v4LXLr+DCs2dQFAQlYaNei50qu6cNKfkNKw8yPRxzdiZqe0YkopPhNRXlIz8IEisawEEC3hTIOSdS7X/g71mB2O9He2FJ1iJj58ZJsACLU6BrL51xFu0ZaAMQS0lRdNoGRKOL9ieG47/O6kVBG3QP6wCyRSo+uflDPD2IYjqKao0oTxxpfwojKfNKWRQlYenYDBaWZ3Dx2ZMYjsYYDccYjyoYY5xSETzVgXb3nIlZQvfc3yHu3m95RB7QcLP1l8TiUuF1SlNph71jHYfQ4bvLoIk2ZEb54+l7lPPk2ORwxxG0ycuePNcG4EGWGryruZ0UR1G0+BRGGg+oxJE6FR/KAwmx1AmAkP4FPuLRTFPhlL64c41hjMc1tjf3cPPGOj7++Ao++OBjfPzZNayu72J/NFTW2r7O5t6a7c5cP1EW3xhj1m7evPm4i0cdmh4HAMh1Z/68Jv23u0N7wrDKdZZhcXGAl165iNdffx6nzh5Db6YDrQElE3UCvNZQOWF5eR6nTx7HwtwADMZIZ9igDKujCsN1YFgyFnLCwnwfJwddzFuDkuugoEV3cSCWNEs9WXUU7LD+sN9TbyyOxIyVAgA/Wdwhg7hhHsQfkCBMDhq0n4ptoBqu4uTINEokXTiLkC4essb1jNo6SXSzcVdF17twLACANNOcF1UheiJ59rB6mk8iGEpJ3Dcn+5mJFhAzJEpiF04YkoSxJeIh+D3E/rGEVqZD5L3hXfck5DPzIIUAaMASjCHcvrmB99//GO+++0eAFF6//Cqef+EiZud7ANUe39gAaprMZcp74tZRFtuSKyGtlIpzgOFMvX5Dlb3visyPEJQCdnuScM6mNpkxoLjTFGYBA5pDhgEXAUDihqpCFH14D43RdEfcTlm05FCKXIXRU3y+xiPL3PMvM5hagzkqbivJT3NbJz4bHeRqITz8rnTweuL2IpTTEnCrNFB2GUWnAGY73mkxOtSmFypIBc9EpDcmpQkHp3Vbxt/651XBifLulPaF7gYApmChBqSkNrSb3kYAeq3rJFjhrveVlya+VxzfTwOQ+T1S4ecOAMgI6cDJCOzTsactmHibez1Pu5sMGP/yrCGMXjJ49bXn8Oylc/i7v///8e77n+L26jZGo4pur26Vs+ePv110y/dVr/chHn2iqAemRw0ACBj069qc5yx/qTK2CzD6/RLnLpzA6288j9Onl9CbKaAzx+STKucJub3BotTo9jKUXQXSFYzSGCnGlq2xaiqsWobRCrrMUZYZygzIjIXm5nLXQaghetiHiS8Lmf2Cl/6Izmr96VELDRbKxkISlM9xMvtZS+nJgRFGpNmc8X4/L6DoBPum5wXg6p+NZR+QozC2IkR5CpNM2+Mpx+zkMaSFb6LAtsSxz+E5vPgInEC2PyRczXmTp5aBsL8cPiNKlgA0ZGhTgyelZyRCdTIOHVBuH5ABYg2GgrXAndvbeOc3H+Dff/0e7qxu4plnLuGtn/4YJ04vI8v9GJKEQnIca6d3tG8SeyavJD0Gp62raOJI2uMJVCj7tQKO0uxrCOOXOqnGe4tjlXjWiwAPgDR5GigGDKOxJiQnhvetSZ0zJ0RfgkUEgYSIAo7xAlHYCBnf0eDaGxqyAAxFmNeAKwF8TNiXptDhHDUD8PVrX1Zw+B7wTnPySXrZaCX8qxsvRSZDC9VNkIvqUXIdAzQ1amQaHQx0Qu844W7JaXFGYMq6mbyNPJuUAw5AsHm3hM2kSofczQYB7YaoPSYU+kyIvkHOt0hiLqyHsuR8GsIMux+x33g0yDaf9ydElmlkxRy6vVdhrUVdGfz29x9hY7MiUwNb2/vHqhG/WGp9AcANAOMHuvkjpkcNAHRZqnlr7HkmOmaZM52DlpYHePbSaZw5u4TuTAGtAUoWOsuiSCcIWRSlRqeboygAqBqVAvaUwp3a4uZ4iG026GYavU6Ofq5ROHYOMVmLppGyhmDuTwUZA85Em1gAUoYcNJKWJp3O9tQULuF8vv3ki4aQbPQlcLfk2gSdw0/6KPhbffBtpOChwfMaayEBFK37HngM8OPaFD5iWLYibTgu0BQlBVMbxb+bgYLTQEpzAQcDDktqoeb30TogYzSFGUropte0Tc3Y2NzFu7/9GP/033+DL774CnMLc/jzX76N5168iMFsN4n5F3NtA+nck9Lwo/gj/uKTTKodHOACZChaASSvtEt9EHridqt8RAlFbUgF73rygjsBAOzEnE3e1SS6TaZb61h7ptPEWeEhmtaZ+LSt39PZdvNbAV1imZOtoYPex/0Igru/W++i2mqyrTGnkEGF8+Oa8NsAnj9NkmQStaENpubopnDvgcTctKVxP9e3wd5dbxWtp2LuYkr98KUhBVHCpj2fW3oR+McU6u79RwBzWLDU7qf717lUcSypQQStCF2tUBazePMnL+Pm7VV8c3MVu7s3YSvG1tZuRw/yc8vzK+eX3pz793feeeeJBACq08kXCOqUMVQSKSpyjeWlOZw5dwLdfgHlM5CBVOK9yh4JxgmiNNDtZOh0MmjtzhuTxS4Ba3WNO6N91LDolCVmOzlmNCG3BoojEo0te6e0aXaphrkxubDFBGM8fTiACWbRkMVxhcRWkvu3HQCofY5c214AaeeTva5GD1MNZdpisK3z2mF1Uy6Jy9h9YgTzbupDEf8y8Qk8IGoOv3vzsdA5e+EWu6C8xk0exDHHcaXwnlXTiSk8E/tRUY1hd+LO+XTUFWFjYx/vvfcJfvUP/4JPPvoC/UEPb/7kdfz8lz/Bysos8lwYvme+Qc1ti/Tp1PZoDldQ/B1HBFF3kf3h5Giz9G0LLfn7EKUC3++fSpyWD++MEQXO38Iww7RiNSaIJvX29qgCUSwn3fIvNQqz5hNz46Mbn5a4T4BDTJGdjD0fXJL5MDQtYVDy7ZSPU0aqYbUJKBjN9NBtYOVB84GdT0F5m0clfKKxsA6YjwnzYGom9XqgseNoPZjkS+37ptZE6atNeK1vIOWBjedrK16TTxn4Asn9HmxCcIJSxd0pjL1iaCKcPL2AV155Fh/+6XN88eV1DCuD8ahS+Xx3ZW5x4bQZ7xUAjmQlwkcOALrdcjDmbHlckyLSKLIMg0EPCwuzcJkvPQL2IWUSJx9nEYMUI8sIvV6BsiwAcgxmrBS2QLhTG2xXYxCA2aKHuUKjR4zMmOChH8QvOdEVzeNTek3JdJoym1Nz0r13x9SE2G/GKyeiQGZYG5hwZKKc7JMjrJfYP06sE1HoHwbLS1JA32JTDifP4e6d7q41IArF7wWNx19NQ7lcpNL933BYRlbyJ3A4JrHByTC0ntGnRg37nt7r3vORNs9mS6jGFqu3t/HBe5/gv/yXf8AfPvwYs3MzeOutH+Mv//pnuHjxJLJsBFDtmUo6J+Tve+Q1JgFKk3DyQC0l9bIP4Cm9Lvmh5DCoiSfDlLUwzC3fgnQrQUDAt9uyZBIA19yvbm9yTFAyMZK3jLCFBJeY2+9OHHz/qds934bEo/9wNBVENCZeau+abvmZvLgp4qbfrw0q7tau8mvJhPf1wCS8+xDnNWd+i7ce4NgxMZ409c+k1Yf68mPLyTBJarcyz3D6zArOnjsOrQ2kmFxZ5nOD/mD52vrtDg7PiB8rPVIAcOrUKaVU1q2tnrEVAHLOM3mhUBQ6eLAKWovmVMnsVjuGT0CeZ+h0ShS58zy3SmFMOe6MLe6MDcaWUGbAfJFhVhM6sNA27pvJPleTrR3unbi9JJmswfUJCD1NEWa6ENvMevoxCQ1sL105g+AVh+Raac2geRy+V3f/PPmE7t94XogpngBAk2OW4owISGQJGsQSSRzzCSAuUwr3iT1JcyY0dCUBPXxXsRl65uYYN7rsoj8cxzIG2NuscPPGHXzw/kf4r7/6Z7zzzrs4duo43v7pm/iLv3gbzz9/DjoTh0EWP6Sw9353jfFuFDXxNP2YRKm4IA2pctfe9U5Co+BiCGzgTsqfkSQjSyYXsw1gitPv75MOuoT9Gm7d9p5EQFNoJy+eQ7sU/z5y7PSo0rSB8jz3wO8P086jEbJHkQ58UnKWgNlBFwuLA2RaQdEY1gJK626m9Wxd1yWeRAAAAER5RtAFg8h5JKsQ7xpZuEvOQz7jXjMO1YJIoVOW6OQlcqVBrGCgMLSEtf0xNkcGTAqzirCUafRAyNgJZ+UZhbDOpghtM5EmuxL9wynl/m9ql1EF2mKIIEFdbWqbOwFm7cLbArJs9SkxCnC8DCJEdeM2D58pTtZcbIvdqOEzJJFG8h0pv7/uNTJWE0xegSbuo1yyhiSnUIow2tp/BI0B+YeMj7LhI2q3q3pmasZoZLG1OcRnn1zF73/7B/zpDx/h6pWvcezYCn72s7fw57/8CZ65dAplh0CoEefHo2N8ygMAl9y25TCVaB8p6272yp+R/ArbC2FMDNpWJpr4cK+JFIX8oegwsoPSmcOS1ypwTgG8BpJwqK0Vf5/o2/X9/kHnZEjd/Tump+c/2L76943ScRa43fzsIGmmFHKloYmC+qqVzlSmOkPmAkd0oj5SAGCMIV3kiqzSzvnOMyBLgFWwhrzzB0H2f1TQXnxIDSlAA0Xeh1YFrFFgSxhbhT1mbO/UGO1ZFKyxkGvMc4bSEGAAVy6oOe53NVNNuPO7kyWTnZxCE1MhPXvyOCe/GYkx0YdSHcp05hsQvS8w/hTHHGDFSzBD4wBN+671vdtzT9hGi/FY/xyE6JTXXCLkg/WSMSUBZU6gS755habG3/D/9mYGn6YjyKiUrbnuSfscd5KkPWNRjSsMhzU2N3Zx49oqPv/8Kj7842e4cuVr7GztYH5hFm+9fRk/+8WbeOa5MxjMldDK+6M8tkieVN9tHxeKWnwkCatLR1u58WL4MZGtmZiDvYE3KbErEELM9SQdYtJOVf9pSq/TC2z4s3lWS+Bw2wpwP7aGo0CPVh5MjWRMbzk1Lu9IyqjvjKaOhughFA+I4uGyOAICspVWSqss03WdHdTcd02P3AKgmBWRUhLDbAxhPDTY3RyiqnK3NyvaCgOubqZD/yADVjWyAtjr1VjP97G/Y2CIsEcK34wt1jf3MdyvkGtCMVPCYhdbygJmjMKY5E156UQupJC8xaHNkEIGKkqfIS1x0nLCS+igNzwNAEQBxo3Qm7u3gMDMRSi6nQFh2QdlkmsqznIgfY7UCh3DxeIJPv1Mw8gQf0uKU6SW7AOIgn9BGqYHuDCi+CRi9E4EEDlNWHYu0zsFECnHGKjZgtnAGIO6rjAcjrF2Zxvrazu4ceMWPv/sKr66cg3rG+vodUucu3ASP7r8Cn7xi5/i3IUVdPq5c1JVzi++DQwf3PQfaQIsOlU9AqkkRA9wzw92iXvI2pA18SBS5OxgDVjlkVH63g8U8sRThcm9qLXrkj4hUofYyRE8qCcqMlp/HbeQcxNIPKUI8al1TIgPOH4/7T1hREl2lLYgaEw7V5ZW61zXNT25AEDrDGSJwC5n9XhkcevmBv70h8+QlcoVL0EqbDTIuvSYzlRpoErgxte3Mej1oDLlAQDh2rjClb0am2OLMlNAv4OqX+BLVOiYMTLry9MyAFaOEZIwc4A4Nee7t6f8/I4MX/nEG5GJevY/ocnIdgPQ1OrT81zzUYNtxMsn3ryhaEWYbmmfk7b9eTGn9vQlatoHEmuCJTQsEX5bK2qCDTw0XYNjuSlRsg0QnfbuSSxpS8jfwVc09Mk9UlJBIkUtlpIMaYCFZYsKBsYaVHWN4XCEna1dXPv6JtbWNrGxvo3trV0UZY4TJ5fw0suX8MYbr+BHb7yMEyeWoLPaa8nuHu3Usg9D+ANNnsEUPamDr7jPfBYmDFxeCbbsMjvaaCp3ZzTtL7LdRtJqOM+l3zVihWqBG6iUykQAACAASURBVPh7u2ic+zD1I7EWtQ82nluc+g4Q+EnCLvGHkB/ZHpmMU+Cpc//JIkJ0gk2p7WjYtpgcZtSeDLP/3ehgsJycAz9nlSbSSlttj+zAPWIAcBxe9BDAMMZgb8/gs8+u4vbtW1CZ9dXL5HynjjieywjhQhnQ6eTIlNMeawWMiLANYJsz1KyQEfCJAmYUo+ARNFdQzFBh7P12AjywABD2MBNpTYngY7Je4Drh4gqctDJqUcpwUwAwyVAFVrQBgHiVxwIpDEsUwIgz9voqaZyGPCGclwpvSymQicemkVxrwbGN0D8BRYnUOIhC+6oBAIJpf+o1aQIk1xdFIvgsjLIICZem2jTjuBBrbx1hZzmCCWGezAxjDcbjEfb2RyjyEr3uDM5eOIVLly7gRz96CS+8cBGnzqxgdq4HrWuvhft4f47vSB42zRZ3WDBw0PCJFi4Jbgh+2yRhNiLEGRbMDuBwavQ4gCiUlXYdSFO9tvvWFgntzxMP8sCSdqrKdIirmo6LFJCPhHgCzTjyJ4O4+U8DcDcT7bTf7tSW8KRDqDa5oW0qcULTRirAVnIJ3zM+dNamx06PGADcBLAMhMShTnOxhlFVDG3ZCyk3pBYM6+OkXLisD98yBGMtNIkfPqNWjlV2YIObF4gwIoOKKyiWetJJ9q6wBsSsWft+iobvtaaG+dJXimLJqd2cCE6Ap8tMXn+MFgiJdn12wMSIiZAxkJNjMC1rgPQMoCRtKFiqj8f+tI106bFpJK3K1ohLTSzZZCzIGqhGaweR5HJXwYM/fMNGjANTmvH341Rz9HNFyd/TyL+L4DQgliQLRRakLTJFKHKFvNAoOgUGszM43evgxMljOH36FC5cOItLly7i2LEFzPQ7KEoNrS1CQba0CM1E+N2DURC01Pws2dPS9sWpMgvzW57Zwiq/TRA8/CZvFACCH3wlmyfRXBNOd2UFkguYfFInB4ClV2kK1gcVs7IqDn3+hPUAEYCxTbJ5Phiw+D6TpLuO818sAJKsyp0FbzlKqQlcp+VleEpC0+Z7Y1qSBQVlNg2CJrLWHibO8zuhx1ALwLBDQwylgCLPsHJsEWfPnkReACHTEzOMdfHH7KybYOu8lctOgZmZPnIt/pXW7537fE8J33TxBC5sKngQU0TFDAZZxtgYxLK5foebm2xRcknF9KlNisqUaCYk4ixhcFJyhaNVIBX2ki0vHDtAgwnaofC5tKeHEdD3JlJenxZnFnZFeQ7DEqTnTnCI1UIwjGmOHUd7R/TW92NAQMzRL8lvkmdL0Qwx2oyLYKEUI88J/U4HvW6OTr9AZ6aHmZkuBnMDLK8sYnFpHgsLs5ifn0WZKyjt+yTviCjpW9wHd7f3cO9h+ADIbYDEApPw7WRGNSgR/NFxz7cjP1IfgSI0dQAAMcGJAI8GHiDEqnOT6OJugBJAyzrS/jZZRxONJOBTTgi3b0dEiJNnYruQnAltvPY9pql1CQJRVPwbuTTcODJxBEdovl7Xtv9I8T4PPG7TuvkDeQcAJkCv8GHH1+WktgWGQCBlrT6yqOoxhAFSgJ5KA91ujrPnTuCtt15H2VVgJQAAsMyw1mns1jIsG2htMT83i2PHl1EWuTcRW2kbsmMszFIyP4lm7OLAE8c5ADAWY1MnAIB8fvLUyz4mk4z74e2Hc7/CxCAEEBHJJ7JJAUDgak6AMaem/dTbPJEIcMJZ8UReNTSZ5gN4qqfPQUn/2II4wCDEs5oXhjz85IWO11wti/0ldSTj0OOGwkYExRoRSrnnUKSCBQXpYgsxcelYOUClFCPLCb2yRKeToyxzFN0S3V4HnU6BsiyR5xlU5tuB8ZnyWk9IClIuOu6fU3gf34qSSdIe0aa2IXMlAQGpg0nD61OgEof32PQJoJCkJNSdaMxLEaRAtCulc/VBKH2au/DBCVCbiHbGgYlqmmP15Gj+EPDjIzsAAlsBwQQ2CkzGZYdWPoetRH6kPIToHiDjfujhKCJHk2IRKyvphxkgy6m0QXMMiABS/ORuAQRil0vZoiiBxaU+LjxzHJ2+BitXujXoVsncYTLIc8Li0izOnz+NXq906UzFYazhIe1UKSnMIQxOsc+ZnmrdjICMpTyuVFGLefZi5ruYBKj1UNSa6ql8D5Qy0LsAAJ+O1h2TVKZewPrZxnLTcC8RWqrR3kF00PKcdGxJx8qb7zkatcJZkhshSbcs17oxbcqqlFEHABClLVSSNZE8cws+AOQc0myQRdwKA0+Emd+7JzifgoknZiAkHRYnwtbrtRKqEJBNWhRmSpv3Q/dIo9vsK4NUCgLcNg374iTJiR7AJREEifiXVMDuKQRUtZ8jXXyTz/egFo9Jt9FI6cyNQyuqKeI8av24i+lwSfR+qMQEGLcFUNWMalxjPHI/dVWDySDLgLKTORBc5shyncx1GeeHJbBjZsEfJgiIxHAKTpDsRJAy5Rx4jwIpBW6HqxwhejwAIIwSA1SDVAWoymn/UuDCM9o4Ut6UTwBjD6T2oBW7xDeCfr2LmYQIRYWZ4qRW0mZkus50aLxgtz4s0CWNcSLIlxDy7SlOGXbzXTJiTQElChQ1Bd9B5E4R734VueAB104cZppgynfD4Mqb2Cfjx5tOgKEtDrg3+kUkYCH1Pm9cRxS3XSTdI8k9nIubArkSqoGjpxaQ8IDBN0Puq/w7F4sKqwTUkUVaQS7sxCXShaDhtjjukUOQDxZaj5pSawSIHCOhtFiSn8fhimQtyNoghpQ+doA4zYtAB8zPtFQvovo9dU7y9EnWPnHqOdMOxvoOU1v1gEx8FUh5ZDAFlEx7c0eWA9+T0mdJlCRWYKtRVRrbW3u4fWsdt2+tY31tExsbO9jb2wWoRq+XY25ugIXFeRw/voyllQUMBl2XiVW7efMwx6aVX/J7TQ3LSBJqPU0HaFp4219nR3b6PS4LQJNlsYRXEaCm73m7sXdVsrRHWg7we+98yP6WL+biHQRTc32c3q0fsgCM15RsMmmlpr0NZjXrNWwVWkwFh0d7osIk4VqRL00TyfGYaLqyd3AYsRM0JhKNmZJ/kzFs3VecJaMRgZt9SfvMSFR0bhoe5IoJy0GzlxFUuRBQ5xITmVgw63rOH9Mqp4F/ro/ueTn53jtVkvQVjevcFoJGc48uPi2l4adTwECcLeTD4VptPOxN5oBgk9DU6MEH97b8nGWxlKVzOj6bBoetm9Rx1VkIdBISSo0oAQty4EjmNbsfqTzX2NsPcCRlkqKOt8dGT8LmpNYAH6jGJ31P3wGJk2m71XTWxLJZR5b7HoqaY8yswEyoKsbW5h5u3tjCn97/DB+89ydcvXIdW+vbGO2PwaaGZYMsVyi7BfozXZy7eAavvvIinn/xGZw6t4LF5R4ojxxN/I4ffGqbe5/yPaUJownE+ESBp036bzEs3zvLy3dJjwkA+MFhYV6cmDDTLYBk+NKiNpD9/FgvPlbyS9sIU7l170Rwe1NyPJ6GD8UrgrszNXqV/E3JtU0Nqa2fTV7bOtaYXQxxKoxx7TK54rSD77P4LjQFJjA5BmnvJtFqHANKDyTX2ubJXms/6A7Na8RnIz0z6TQBCGGfHojJqfIeGg2nOQLF81YjtdIQqURIpgPUMr6HG03rf/qpnY3gIRJN9ApyZNIDnuNQyXlEIB/7LY/jrk0BnIuqYONPSO8TLElSzVHyMEi2wda8DTeJ/hfT5l9YIS1FaqqWf6ClIM6JAEzDj2hjNPF2Aj74Himj996LJ5cFdQzc/GYDH3zwBX7zb3/Alx99hdtXb2BvbQs0rJAbQPuETxUxRpnCeq6xduUWbnx6Ax//8Qu8+sZzePsXlzG33EVRElRjK2xaP+4x+4+0mHs4lKbTAkRqSaAz0Jyr4ZQjTY8JAFivtbtJGUr9yvikm7mKGtqBuxo+hanE+3qtvcFb0nA8QLSYyAS8pcCfO8HmWxpuqjuE7eB2EvsJDnMfx7jloBUUWdH2UrYqWmzM9Jd8E7gdte7RiP31wlR0wRiS117s3OKe7d+NAUJbMwy3SrALN86PD9w+1AyDa/Wr0afpjDL1QWi9wSlvvN3jKUdTZsjtcWnPh4dE3kpCQfqn+QAUXNhburevQNBg9u9/Cv5z4YTs3Utl7fgfjyY4MfGId70lDuGJcfNhEvSlYyzYQMUvGqCE2xcnn4Of3wEIQbakSAS//xGIEuadvCdOi2d/34kA1rBG4c7tTbz3+8/wj7/6NX7/zkcYrm6hs7uHubrCIgiLqkBHK4AYY2uwPaqxtl9he2eEL9f3cOP6HXxzaxXIMlx+83kcPzmLslSQUsVpdEC49xNIsr5lNsY4I/l8kL22wdf9zD6a9OgBgISkEjcZT8gwFhnYhCbs/zVOLfHfRTNLIw8+DhIPjqvEWupyppxIzWNoMqpg1Jy6Bg6rykw5Jp6kjfvK39o5a3kB5Bib1/SpeU3M0XaP+05o9AdfFyFIeqTd20MSxVd312sJPgfBYe6Swrz03Dh+QAqq7tJi+PKApZyEy0mb35ohTkFEE+Fs/peMC5PyQtqzHd+GSz6lwqVRUJPzXfFrjJlgmGEaglru54SLtMm+bkdqJ4vJkKatpaSqYRAg0YnW3SaxljXGwRtSPVtQE2PrrIXBtscxI6CF901hV5pV1imRBnHbHPt9J2fl2d+t8MF7n+NXf/9r/OZf3sfW6h7mxwZnQbhU5Hi2k+Nc2Uc/dyByrza4Pazw2XCMK8Mxrm6Psbq3hvd3htgfj8HM+OnbL+PYyVlkhUqAbvPeTzK11ZHU8U8Bd5lmAqWqg074zunRAwATnePcCm0VIYmqjOeuMYGO/DCTTxAUJKDo91N83tv7uXdl/3elpi55WJo2G77tAqIDtKKjQNz6nX7TBFWHaeWe59/txEMO/aN4Q/dHXmh7cvhWQCl7UBu1c6ehi+bvFhOzBawLm7XGOrea1LzvnQZhMpgqw3ikYTVgWKOqFGylwEbD1ArVmDAeuWRYtSX3fa3BRoNNsg6DNSCxSATIwUh/mZacp+S8kPmSPcDyZ1jjkoRNI77Lz/TzW5sCLex/ZOhQy9rNF7aEzz+7hv/2X/8N7/76fVS3t7C4Z/BCkePtuVm8udDHC3NdnCw7zu2MgNoyNqoan+8O8cfVTfx6Yxd/rAxubezio999hG63xGDQRX/wEubmOmBt/a4bx7nYYNSPyPL1g6WjyrcdPZYtADttpU5ZnUHbSrRNEfIWziNcMQDlK5WFbzyDmXDmSu2gNLn4p0xkuecDTfEgpL06EzScye7cD8XsXkeT4l7zxDeP5H4uZ8JkmGG8p4y5aRrf6P6X46NhdpNtcsiYkPbRa9PWwowr1KMxWDGq0RgwzqfGVBbj/SH2d3ahNYIZ181BV0Dry89vox4CWjup8NWV29hc3cfeVo21W3v49ONr4FGNTqFhLOHK1dvYWN3F3voIlXFAgqZaZ8QfIQHtYStBcjpEp05J9CS2BSdXYnvWWOxt7bk6B+4CZylLvNSkXkIomuSND+S/l7Da9ghLyuujyY69xUpsLgELMuCzkFqrMNoD/u1ff49P//glqrVdLA5rPKMZ/9vxBfxseQbnO4Qe1Sh4CDJu7HIAeUYYzBV4pn8Mx/o76N5ew292dvHNNuOD332EM2eP4/jJRfRfvoiMFMRCywdXdHpKAMQQR/Hj1LOInuQtgEBiVvQhdvAsgNDY104MmA3rrOMFkvYnFdNisKbGZ8d0RBjI50h3eyOHZfl301UCu0w1ofuQJQnevq8+3S8dNA7f5n6PdrY/QM88T73faNxvO+ZNr/lUgCaWEYbf07bJN6kgMKirClvrG269aMbu9i5sVQHWoh4Nsbm2BkXGJXxR0XGPucLajRw76zsYzHShiEGksLG1hytfX8fG1g42V3ewt76DpYUZdPIMDIX1rV1c+epr7O5bWFY+3bAX3o3EDt4eYaMzoPVaPUH5508y0QkA8Fo/k9umcFczYBn1uPYrmyFhjM334Pui4NKFEvsiEjE5S3rB91JXTfQI9tp/NWLcuLaBP733KdauraLcr3FOa/zV0gB/cXweF0tGzw5B9dhblzzwIkJBGrnW6Bcd/GRlFkNbY3M4xNbY4s6dHfzxvY/x/IvncOHiWcwMSgB1VGa+lwP4cCnlZ21DbFqXhSFxEPGzK+Z1dGHUIwcAzExg56fM4cclInFcWUS+/zfMO0GizbrokyM5aah3zJ6CJvB4rX/NnnICcH64lI7yo6egKU99oSJ0Enq83WtSct+4Bjw8pWBcdz9h7ru02XmuoJQFuMLWxjr2h7uAAsbDMbiuQMywxmBvp0I93nP7/Qo+wsPCcg1lgRvXbkITXFpnpVAzMBrXqEyNLWxh7Zs7KLRG5jPGVYYxHI9R1wTnpyMdbYJRsQyLT0LYCpCtOn9C+N4fV3Lc/21lZMQZkQBNDNKELCNonQxj6jzqwZNiC8VJGmeWyIgk9we+uylwb0qjWoR8v9lZNveHY3z80Ve4cXUV9dY+li3juW6JvzyxhIs9jZ7ZA5l9wBi4pFVpMjEDqjV0AZwoenh9fgbXd/fx6a0tbNeEG1dv4rOPv8JPfrqD/kwZckeEnjw1+Qdqz6Pgs9IYoqCmTrFFHS16LE6AZIiY2slH5IOUW3XauqRdDeZB0ZCACac/YZ9B/AcVIH7NU7wE0rt/G5q0PrfMpGLKe4CbPa5p8+0Xt1yvJ448SCuHOfHA8UwlQ4sO5Yj4CMmlOfZ9kXlN8Kl52S8DCk6n3U6OwWwXM/0Co5FBNdzBaBjD/DRlQAaXC8FajIZDZ3YnQZyidQOj/ZFzivOOfKw0FDlhb9liVBmMLTmNnt1Fzp9Po5F6iAg2FIyKxCmI98KDbBD9yWvx6zxVLi3guxIsfVopaGXR7ReYm+uj1y3ifRrLm0FsXNXP4CgoIKWZe+DIJmNt86zwMSY3s5awszPG7377ITZXt5ENaxxXhJdme3hlrofS7AD1EGCDGJqZmhH8uFUj5EQ42y1weXkB/3hrE2ussLe+j2tXbuH6tVs4dWYRSj3V/g8iJ52aWr/4o5G3lCX+J0QUM6UfRXocWwAEUtRMUZpWxJum30dBKt96Hukrlh1dLP+UnlKDgtncC29CALlyQmAcHBnJYLaH8xeO4/kXzmL11gbGtW1AWVemWszrnhkp3TCBs4XXjGO9jDR9tjj1gQHlazhLciZmhuKm30nw45eUGtQ0iQbnMcXQVqH24b+HkyQe2TE7Hw9tcOLUPJ59/hzmFgaJdi+Z8DzIIRdSfKSV1Da7ukdfwxaI53/WWGxv7eC99/6A3fUdDMYVTg76uDA3gCILmLHT/MO92mPujdOWgWqMmbLAqV4HizpDXjN2RxYbd7Zw49ptsH0J363J7GhTtERFq5dUmpWEVhSc2QGAwKyPbMLqxwAAhIlQa045jb+1w9L67MJSLFPIzBdL/LVu09r7e0pP6bsmCd0EAZZSq5bTxFWmQNoJMGtq7O/toTZzyLVC0Slw9sJJZJ23sLW+g7qu/daZk76KNZhrSKZDSeTTTo5P1gMAL6kVpdEHcRFlfn1KvgBmRsZZuC6UHkYTpovMB5KyV4qhrIIhm1jg0qwW8e7hmC/65DJCKpCqMbfUx8rKAsoyc5yCgfGoQj2sgu9AnmfO9+FIU8rrDlOsy2V9FN5prcXe3h6ufnUVvD9Glw0WNGG5KKDY+NKpMpptnpp0wZtcFBmUOsdSr4dyZ4iMCdWoxs7WLqwlRKfEpyBggghAw2ktCZlNrIyycc0M0vqJLQd8HDFLX1PXd5/bFoD2d96P+C7zUBxV7+L//5Se0ndGE6lCPANRGujPdFCUGZQiDEdjfHX1GpZOLKE/U0JnCr2ZHs6dP43qZO3D4xRAOhSnYjYhxTKAJCMgySZayLgtmjMltTHSLmnX2Vh8hxkZqwQAxNoYbbRNVvbc5TsLsIZVNnl+Tjzx/dpmL67IVeNkOKCiQQAZ5KX246NgLWM8Mli9tYY7q+vIVAaDGrPzA3Q6nW//oo4ikQFDwTJg6hr7e0MUxrlRlwou2Q9wMIOM6qr/zM4sBFcxs5tnyDxeGI8Ndnb2UVUGeQEo3Sz+9ZSfOpque7ZWOYdfxMxPdjVArh08OpzVnlp/H5BpqbnNfxcY8ZSe0ndHMQogtWwpV5UvJywtz2FubgZFnmNvd4gPP/wMiytLOHFqGf2ZLrQmEGXI8wzI4W3vbm+bJLFWAgCiBogEAMhess8dQNEKIPH4hGauDqk3oMSTn20Iv4vbd86JgZj8PaSAkTfLs/ZWD7HYuUqEISiQHADIWLkCP5ACUj7dNzuzPltGVVuYscGtmxv48vNruHnjDrKsQCcnHDu2gpl+DylTOHp84LCav6OwRZP4ViilUJYdQO3BgFABqNoOFEheoty34TATt3fcuNawcBbWcc3YG9bY3t5H3imRK4T3mUYDPrkOgc13EojTVRcOeYuMBSyTUvrJBQDO+ihFRcKxA1bpNH+A5rep/fGp0H9KR594ym+G1oRjx5dx+sxJzM1/iW9u7uDKl19jZtDH+topLCzOoygzv4fuiEAg9gBAnPOTKmVePicKoRPO7k/HkBhSplREudgDJFYfkGTbiqRCn9+m8CsuFj8haCIQZwgmfoLfr1dgNtKNZunUxrFYZiuYqGV7wDNXYxl7m3v48otr+PyTK9jc3EG328W5C2dw+vQJ9Pud0P+k+aNDDcZ1H5eRy5CoFKHT6eDEiRWsbl7HeKSwaQzWqzFYdVz6dKmTbeWGia4qQksRQApMCpWx2BztowKjAmBYobbAnfUt9GcXobSCVkdsHL9T8nMfMVWykJQ2l+qo7NeV81uzBFRHdhgfMQC4CWDBD4sUhIliWzSY9uik40utb+RqZ6ZMzjuyQ/yUnhLQNh4qRVhamsUbP34FV766ifWNP2A8GuFPH/wJV7/6Cv2ZHoq8cG4wos2z9w0ngtbax767FWFhpmS8iIwoRNIohmKCyjSUUlAs/gHGBeey08GbNczYFwaKgl+sBxo+3XAIEaSG0+GUR596LAIZl9wLcOWrFRNqY7G5sYvV22sY7u+jKDXOnF3B//Gf/xrnz59AUSoA9YO9liNMom1qrTGYncHrl1/Gv36zif29XdwYj3FlawtvL3Wh8txVfzRtH6oW+CQN6BxjKGyMx7g9GmGYdVErhbyTo9PpYGtrC7u7HeRFFzrT0hF/vfPReDKZrfehCR4ssTaAAvnAG+tTA4uya0EMa4gOb/55zPR4EgEx2uzAk1/swfu5cYnXJtA6yNFkmTR2ZEf4KT3hFIVxKvSUAsquxmuvv4CtzX2YEfDZp1extzfEcHcPw929RtGf0ESykFyT0VvG7aenhuAItqVQkIVzshPrgfJFqcha3573uyEg6Ox+3TV2/sWa5zs1KRMmpb4cSeXJQdhA7uuiJJVzTmPG3FwPp88s46c/ew1/+VdvYXm5D62n3f+HQQwAitGdLfH6Gy/jg3c+wM2NNVwbjvHHjS18vTOHs50CncyZ9UPZqzDtkgmjNGpd4sbQ4v31Hayywh5p6E6OuYUB5hdmMRpV2NraRa+foyi1nw8G2gPDH+xA35MitG7WnG2m+Io+MBbWMjOx0cwVHsQE9BjokQMAQy5VR4ocwx4Jy7ByYFD3tDlJ1TOKMdPS6IPE2z+lp/SoiA5IAUZi6laE5ZVZ/PTt19DrzeDdd/6Ez7+8gp3tXYxGFYyp3cpgZ/MiCkZIny43CZONyjmASUWNfBSNZY6RAB5QAACsVNOULIQElgieVFNPnkMy+JGyE4I8deIVapdTTY8JOc0qeQg4HUvpAoNBD2fOHsdLL1/Emz99BafOLKEo3ZaDhFJ+v4mTf6PnACug2yvwymuXcPL8Mu7cvoWN2xU+2Rvhn67dxt+cPoETRRdFrgAag6yJ+6zeUsPQMFkHtyrCe2vb+M3qFtYpw74mzC3MYuX4EmZnezDWYGdnF6NxD33OpyO0J4SmPjY1ZY4T9pR+7VeoBbOxxtTGWl0f1Nx3TY/eAsChkC2kcplL6Su/0738OEYEhFDf+FUKIGxzz4+mbSY8paf0HdPEPlXKB2oUhcbpM0sYDGZw7uwxfH31OjY3t7G/P0Rtat+Ey+wWAIAUBaJE/2DEtpM9+nh/H0IYFETyGQMR1fJGTYeo64hYIm/qlOhG4wW89jF6nJTjFgtdmn9f2UQJ8Mc1N5Y2DBhZC8kTCJkuMT83wMlTyzh9ZgUnTy+jzAEcXevqfVNaGCmCGQbIIi81Tp9dwqs/fh63bt3Bzd0RrmwN8f/d3kBZzuCtpVmcKrvo5hmUHcNt03hrjtKokeNOTfjNnW38t1tbeH+vwmZRgkuNU2eO4czZ4+j0cjAMhqMhRqMxrO1CKxFp1JgZTwlxIKaasBjWGrbGGmPMkZ2kjxQAGGMUs8qYlHYeEc5ZRXbylU/3K0Ag7HUG40qLePJoa5frKT2lI0MhhM5/jjOXo1BVQF4wFpdLLC5dwEsvn8Vof4yqqlylP/HGh6S6jSF+zZulZUqjpq1CnR7VcA6MCcrdv1KKSBwDJcagXZ43TWpkiWHJ59xj7yfghY5OHlrSFSmfk0DuyhSBAvxnw+xyEqT3BCFXGTqdEkWRIcsIpF32P/J9P6gy+/eLOPmRWHz3xrUm5P0cb//ZZdz6Zh17G7tYG97Ee7tj4Jt17FcWl+d7ONnNMKtyFFoDcA5+OxXjztDg450hfnVjHf++s4/rWY79MsfiiSU8+8IFnD53DFkOsDKoaoOqHsMYgzzL3NzxPXwq/CcplvJuHWeGYUNZG9EeIXqUAECNyrKYyYqestSNLIYds+A42bnFflJ/YUoHN1V2EP8WZpLSkR3xp/RE0DRg2hBToVCO+4Z8wH5REvI8B5CHMDgtmjghhOhN0z4k+a2L5XdfKOu3IsIxWV+xAReDb1w/0hK/yXZBtCN4C4QX9EzkNXv4dWwjcAiW/AgmJkLckgyIAGCZtYr28wAAIABJREFUndaZWDSIyOUaAIPINM2wwA/KCuAoPp1wQgcAa1x6/jx+/osfY3tjB7/dHWH71g7+uD/G+PptfLVR4IVBF+dmSsyWJRQRtqoa13b38cnGHj7dHeKjmnE9y7DfK9FfHODVyy/jmefPY2a2C6gaIIuaDYytwdaAWU+E/k3d1np0g/H9oHQA2K0kw0SV4ZJZzwEoABw5X4CHCQA0gPLMmTOdfn+lY0zVHRlzGtAvkqIV602MwoJIOdMWw3p7v0UwUyIx9pMv+UuC8ykwwqf0lI4ytfWCNFuYYpe0x2/RwoEAcnvxOmrJRBw9j8kJ3LCIZINWPnP0CwiZ8P02fnos+NyET3I3xDUJArECSQbD1DrHaJj7ZbtZAICzRrhywCzbCv5YG8zDnyM+DMo/szuFk/v6a1OHQ5uM8Q+CHzTDxQUcCQQjAnodhddefRbjYQVYwru/+RDbt3bw0X6Fm/sGvx9uY359C/0sAxNh3zA2K4O12mIbGTY6GrZXYvn4Al569RJeff05LC3PQWUEJuP4sIzx996n4jGRagahMggGCnsjo7e3R8d6M7NvPv/85S0iu1rX2N3cvL6/uro6hAtd+U4BwcMAAHp5ebmndX+ZyJzTuv9sRjiTl91FMrQyHPHz+3vjJWNBTpugRj7y4GTi45S92pN8YQEyYDKRVT2dnE/pe0RioQqg1e+GZWGzK+EBlH62zd9Nh5nWNVOO361DybkN5YWS8r2BPcS9aQdK/HWJqwGQCGyf8o+k7yF9N929i43Sv+TBvx8LsQrI8zNg1ZQ2vsc0TdMOxxgADLRWWFwa4PXLz0NRhrzs4YPffYitm1u4tjvCjapChyvktVOYKiiMM41xlgNliXK2h+OnlnDh0jm8+solLB+bR9HRIFWHOhBZppFlGlorgNShWO0P0T/gsM8S7U8xgoahcGdtW8Gqsz3d/z8H/e7LxoxvjbB7rdtd+uL4mc4XM2V5czQabX/99dejRjOPkb4NACAA+fLy8lLemftRmXVeh8XLtqqfqarRcdJ2pobqjsa2M9yrC5ZwI3+h8rDd8YWEg/GUqURRT3lKT+l7SRQ1urYNm5J5T7JFlgh7uSYceyDywpSd9w2xX3cBcEQhD38oRJDdC2AkS1acFINFgxHT1BNPbSQxBiQ9YG9pkJO4ISAb/IDuASy+pyT4KnwAADCyXOH4sQVkP34JnV4fvZkSX3x2HWu3t7C/tQNUQ9TWwLCFVRp5XqCTF5iZm8XKiWWcPncCZ8+fxLGVeegMAFn/apwmWxYliqKE1hrKK1stC/dTmkLeVu1LOBO2t3aJR7y40O2+kRG/WNvxjmVzu8iLq4POzGd5rj8h2n732LFjX9y6dWsNbovgsdK3AQDF8ePnT/V65S9Go/p/R8WXM0tnad90s/FYaV0DSmFkAV0TlGpWFnPORArRzSiUEsH0KRbTUv0QF/tTelIpBb9eeQ5fxT39h0kuiSAlKXeAqPWLuR1QrFz1TdiJffZml1Qw/TsQoBpnphkHDyK3o5EqAO6owsFq/g9R62zTxLOR84PI8wzLKzP48cwLyEvC2fNf4/q1W9jc2EK1v4uqGsPUBqQzFJ0Oer0e5hcXsHRsGfOLA3R7uYsSIImmcvOPFDDT76NTlL7I0uSbewoG2uQ2vwxLEC25hWWY7Hioh9tjnRN3LNcLqsBp3ctfZcXb43p8tdsd/HO32/vv5ezsb69++ulVAOPH2fMHBQC5E/69v1Gk/x8MRy/p8c5gzkIvgmmJCN2yxCgvcaOy+MJUuGkZdWMyNdWZtmNfY9Klqg8xDrIGHAVG8KgWxFF4tqd0CGpMgESH44kvp17CNHlamn9cMvAhAIUD1kJSAdAdiMA6VBFI2kgzFkgWPwb7cw4C5ckThI7LHn/TuQ8c53Do90Tmr3vc5lEugvZ9H+K9DvtI07ow9VoCoFzK5F5P49Kl0yjKAisnlzAajmHGFcbVGNZYkNIo8gx5XiAvcqhMgzI4p9OQyUGFOVFkGrMzMyjLorFB1ehnOxduo28P/yU9Tp76oNMvurK7pZZZxgwTVpTCMVIo6jFqU2FcW9obj/KdrZ35YUazi2dOnOZMPZMjX3n22Wf/7rPPPvsKjxEEPAgA0KdOnTpZlp3/AEv/92h39NrMyPROW6svFRm9MtPDpUEXM4NZ7BY9vLe+h3+4eht7wxq7uYZi5VG9gpRSBBAtj37Wx0nnz/W+Ayw5zae8qSe3UMVTOlqkPPO0cdvLy8bUEXCCCDCgA3ioa8DNe8nQd7BJjFsCNV0uBhEc+DQd0CFkMan6F4R/bCNoi643Tkix9bH7FErR2zQmkcjn/Zfr4rg0Ht7nBwH8FiEhAhCyHjM0VYiHSRKSaI8oG0mLS7mICAWtGIPZDhaWehjVI+zuADA5rC1hrZ9LKvG7olC8NtleMiBi5JnCYNDBYLaHvMiihaWdkRKAq/LaJj3l2BNCslfGhAyMwlic0IRXZrp4td/FYLSHuh5hs67pm6rClXGlrteV2v1mbWFY6repyPpLc7O9S5fo//3000+/BjB6HN2+bwCwuLjY17p4ox7X/yvG9eVyOB6cA+HHswP6s4UZvDRbYrlUyMsCu7rAeH+E92HQsYwh536/k6L2MX1bEE2WRQ1kOc0G4LYyqXVgSlPt774FtZHw4wIg01DqUeBZ9zvME5rEw2Tuh4Tyj1Dxm9regVXhWydyVM+TE0TD9tnHpsW+pko/NKx3qA15/JkAVrDG+rwABLYWxqfatSrR/K0LDXROfDGUT5FCKHBK1nv3qyDgSbl7sdfypcyvpARrPGMAPNHOoII9ovWikudzKYiT78Kf/spDr0VufaKkb7Gde2mhj339iSJEQJYT5ud7GI3HsKZCPaphjLcShTLOHpk1TauQBFBaK/T6JVaWFtDplNAqwrVHTm2LV3LgwXjqY+aQ7EASsaSpZxTWYk4D54ocr/VLrOgKZVaiKjLcrAw+2Nii36/fwac7O9mwKubV3OA1hdz2evPrzzzzzN9//vnn1zAdZT1Uul8AoLXWx4k6f8Z1/ZNsb3/+ZG3ozYU5/OWxRVye62I5r5FxDcYYGeeY5xp9tsi8BkCsDlcamBGcT1yt8XS1e20IkS+E5EFijZzSXmjhEc6FA812ST8aJz8kuh8w0jQpf/tO3NU4/JDvdT9EDcFAkwcfGcU5Ou2Zv9UoNFBzNDkC0aDrkm0BYIYxHmwzYC27n6rGaFSjri1szTCm9omHDAwD1loYY2GNiHF5FiAjgtIZKFNQWkFpoNAlMp0hUxmyLEdeaOicoBRcSKN2EIR9zn63PUFRHnHj4dy7cqaFZMB86eFk1TfX8RQ0cK+hDM6Kvj0kIcaJFTLM4SNiYQy98NuhShP6MyWWzQCwNTbWdjAeuS0AF1xNrRnjPojhX2tCr1diaWEWiwuzKHINJY5/3uoibyaBWL6hh5N/NU1K+XD4Ypq66BG9N5kW7OSPk1XeZs2MAhazsFghxhlYzOUaelDiYpbhZFdhRVWg9U1U47Ha2R3O7ZedV5ePL/6nbre4urGxsbG2traN+5nQD0D3CwBK5uJ5a/j1vMaphcqqlwqNvz62iMvzPRzTNTDaBbgG5R1QVkDXBpl1CUZkgKQKiCznxjtKZ2hYjSrkMm+MenKJ8MWDBLCkPuEDvn+YdM/pJubN+73uKd0XxSQqUmUeaIPqewK2+6VEok0zQsmx+zeWJiycgYltAABsGbWxMDXD1BbV2GB3d4ThfoXRqMJ4NMJwf4ydnT1sbe5if3eIelyjqmuMqgp1VcNYg9oY2NrAGMS0w34UM6Wgsgwq19CZRpYrFEUHmc5Q5l10uz3Mzs1gZtBBt5uj6OYoOjm6XY1u3+1DuxAzDaUl0JCR+vYwfGnVMGYE+LwComXJYzMLb9H++vuNpor8hB+RgH9Yrba3P5i9yxkx8lxhbraLjAi51tja2MZwf4SqNrCJCZ+9gkRg/E/m3qzJluPI7/x5RC5nq73ujp0Amk01l+6WWtKY6WUexmy+53yGeRwbM82MSeoW1SSbJEDs917ctfY6ay7h8xARmZGn6oJAG2GmAOpWnTyZkbH48ncP94hMwBaWyXTEweEuh8d7jCcF1kgnXsNZdwjgBicu9vz0RifuD+lbbN/3qOhNt9wmT3+ojP3X9COyvCFuoxVGzDmkqcmbmnGzYVRV5DVMixH7uxl382MWolyfXfP5YmnWWb4n9+78L85l/3UyOfjy7OxswY/sBfhBAODhw4eTTMa/qKv2ndG6Lh4Y+Lf7M/72YMaRCcq/WXvlbHIww006B8Zvl4IUhVoUmgEcaCq+/bnj/rxliSjiu4NRGJ7b3LfhO6Z4+/7QtBuGRuKG1ORB1dstvu1Wmjdcv7U3t1K1Dj7Gf3WLE7+vI+xHAUSJ8Rbbtd2+G4FqbzhqVLc+3Gr4bd83eGTroe/wwrz5q61zwP+Msrjx7Q84uzreOjCAw+KBYoN73qAt1K1X9FVVs1qvWM7XrJYblsuK66sVL1+ccnZ6xXw+Z7mYc31+ydnpJaenFyzmK5rGBfZTnAv8qrGvEn5r8tOvK2PEHylsDKpgbc5kMuP4zjHHx7vs7k2Z7IyZ7U44vrPP3XsHTPd2mEzHTKYjdmZjZvmILBdsIZhMvOUZ9wKRlLtA6fcCcQkfatK+wdLA9y23TfqN1LeU577Du3ZLVW+iqe8gwzeWm3VGGx/yzLK7O2E8HnE2Lrm6vGK5WlPXDXWrPQMKZJkhz3Mm45L9w13293YYTfIQHOjPloyRLDeX6m772MeuDEyz7Udv2+sg6Um46c+Ow/Yi8L86EfQ7EMJQ7rzpfTGeTUFdt+UFKE79D85hXeuPa24qqJRClHd3JvyHh3d5Wtecnc+5qFx28vriMMvdLw8Pd/9xNPrwyeeff/4/DQAQGE3yLHtf1s3BrG3l7dzy870pY2mQtoK4ZohBbY4zGY1YajG09GlH/Qln3ALTtp1V2h2CYhCM+vChNnoUSKtR2gGHhNPNNAZXhRXYgSzeVkLBVyDaX9f+0NXeV5Vs0jnwNb9BiSXviEFGt/LVGxVgZLPUVzbc1LUlGbXv6bbc3q++a8vWuLypbbc+m3xhEBwmyJ6h/+WNwOPGMbjbWjqeZtfXl/YjCpkmWDr+m8hHQUl0+8gP2yJJKtrN9nXn3w0Azg91DadC9ebYRTAXvBZRbiu0TUtVN6xWNZt1y/xqxcXFnPPTS87Pr3j16jUnr0+ZX69YLWsW8zXXF2vqTY02Na6paKqaal3T1G3gweCbUw1HA0cF4MFG38ChFSkGREwYa08rDY7rqwXLs4oXX78kKyw2N5AZilHGzv6M2c6U6WzC/v4O9x/e4f7hAfv7Mw6Od9g7nDGZFoyLEUUhZJnfFdF0GxJoctyxV3z97AXq/zMKZ7sYNZ20cRGt3vZMd1IioH5PxcG2xt8D+Mdrt1mm3xeE31RDtv9bBLH+9+HhDpOdgk1Vsdn4+XbOj4+1XvmPypKisJRlQV5kQULf/kIv48IurQpIG77qt5q83bgauuJv2wJa4Xbvi/aw0z/TNyl6PxC/rNxRZ1ePeeOYbl/vUm9vAJg3F78b9+A8Wu9p6X6EFqhE2IhhbTPG0pKhqGv9ltbNhvcmI34ytvz+dMPFesXl+aV59N7d96e7B4+WX1+X/MjBgD8EABjVdirCvQKdzgzysMx4bzai1BZpg4A1BWpzNnbEBTknarkUw8YIDT4gpQX6JJRhieipZ5WtnQPj17ds/pE+lVotGjwN25HH0glyual0SAk6sbNTXb/1+2Zr+mf//P3fXfTGH9tAPB7h0qnEN1QiAyspTdW6gcMgYdjk8sB0Cauy4q1Go6lPYuv1g+duNlFgcHz5jT5vWx5hsrfv7y1+Sd6Zwqj+uT7KfIjK0j1reiAkfb2Djt3sh35HrMFA+W/rrJAZ45zQttDULU3tWC5WXF0uODs75+nTl5xfXHH66oLTk0suz65Yz5fML+asF0vaqvVr+5VDN0reQo4j15aRa3FtS4aQGYsRg5X+BA4VD6/TCJtuXgScA6f4/HEBxfi4AYVGhVaFlhXOCs4IjfE5TVcWTkpLUY7IcktRFuzsTdndnTKejTi6u8edB4ccHe/x4O4d7tzbZ/8gAIJRjs0s1tigb9RvWzvg9n72e76+RTEncynJsy7ORaTLdFFaknfobXUNaSClv+0bPH0n9HPTVXTzvgEtbfsApOel8Ke1QjHKsaUwcjlt43Btf78Vg7WGzPrzJowVb8QmnRBxqCZnUNzSxgGY0a2+poyW0FE3nolyl8HjHeKg5zNN3rP1ZvU5JUNtcDvEkuSd8fbUiOzlQVLNbQImmKORTHqvma/doTTGsBTLqRqeiWVkC0zWsmdzCiugLeJaDgvDI5txpPC4rqXaVBRl+XBUjh40TTEBftQ4gB8CAHJXrXelGO1louXECPtFxmGRYbX1CsBkKIa1ZjxdKV9Ua35zveHb1rAyhlZiGlSwmmNwiUh3ylhPXOFvETAeODg0OEJ7K434Ocxi3ETYX3cYGKQ1eZGldElJHTV4BdqDkptnucf7BwQTvnHb922XsG/qd65acIsja4sxoms2skeAOOGO3mXrmbZvYRR40n8cWPjKsD++r2nQFQzpsD8iVLe+icy9/TS33RtwtHbjGoRt4NbuHdJ/75VVWFzasqRvtnQISFKBtd2zKFa6oB5NjsyNo6zDQLE0PLXzEhHb3i+ApRva3BiPcMHh0XFdOVbrhuvLlVfwFwtevHjNi+evePXyhCdPnjGfr5hfLljPN7SbClu32E1F1ig5wgQhV2Gmwo4IMxFG4ihR8lwYW8soyyisJbPejrTGYI0fW+l4pD+yW0VoW6VVR4MLm58IjVM2LdQtbBpl2To2KCuFRaPMnXKNY7lSXFZRqzAHlrnlZZnTWqGclsz2J0x2J9y/f8iDh3d4+OiYO3cPuXPvgOOjA3Z3p4wmOVkuSCY4AyKpwo+05OfBG/TblEB375ak6euRnh4MfoKcDGnEbNUpTjqec+H3bW7pGFv/5yIVbr9vGwH7f7qdluO5KghqvXcgQ8hywi7r3gsa22XEhCwR3y/XgaUQzY5Dw/btrYCJ94Yx3/bBmNv6FSx00w1qHEEG43yzRC730nUATrT/Pgo0F951s/QeiOgzdsTU3F56pp5AVQlOxp5njQoueA3jEnQvGhRV5+sT74VeW8sphs+rhul8zWutOVHlQyc8kJxRsDByDEe25NgW5I0/iyHLsl1ROWzb6ym3o5m/WPm+AECAQlX3nHMTo2pLq0xyQ5FZcC1qMiqnXKwbvlks+edVy+/Xjn9ZOR63sLIZjYRDfSTsLCY2CH4ZWmBddwNQMIBVnPFulS58AIgnCMZdw1Om9sdYusCYQaQNhtITUWoJAAMwG7Fnr0a8q9TFjwiOIaLvLIAEXHhtkaCH7aLJKWzDL0K9Uat6rjHhPW1sRtKAqHb8ca1BtGkMuBpaENvKyHWWi8e4osP7RVM/SgQBQ2DA4Hv/bNcmzE203z2RqlLXsX3b1SMYSY6avX2k+n6EeJE+oCl+26vlKIRcmDNV58dWI0AU+gNt+/TVtluFkI6C+pEawrJhT/s2SuLibxysq5bl1ZrTVxe8eH7O0yev+Przp5yeXPPy5SsuTs5ZzRdcX18jTjANFCpMRJii7DQwFWFmM2bGspMb7hnLndxwkFmmRijFUWaGcW48AMgNmfVLa5kRrPHxNjKwlEPfjOBaaJ3S4mgC/TWtULVKXcOmdiwbx0od167lonWcNi2v6obzpmWhwqJVVq1SOcOqbpi7lvX5iutnlzirfD3JmO6P2T/a5fjOAfcf3uG9dx/y1jsPuffoiMM7O8z2xmQTi80Eo71wj6clCjf1QefNSphQ0STqP8Jq1814LN0Ob2EwnOuX30QNRi2tajh/OR6nZPqnO3nQn654M+Bt24yQ0JLhtaGZE4Or0xbHXVP9MpJof6BUVw3gcP1ypACStDf2QRyqNpwmCb1nxPOx061xkthf7SqOc9P5KKMcC08O913Yjt7f9oL0syTJ973cortv+DHWZ3C0iGo4Xkr7Meh+UoMukd9EfROBSVriVkAOZwy1zThrDX9a11zVFZ+x4bMM/r5t+Xvd4YNpQW4FkYxZPuKoGFM0VQh+tYUKE2B84zV/4fKDPAANuuecK3EqFsisBZuhqqyd8GK14ncvz/l/Ti/5rBF9KiWvbMGFKaQygDhcAABOdEDaQwXWXxwmAKoX6FsTreH5LjI4fh+3MlU6Sy4KXX+fF92avDttg0qi/KOrXP256tEicIEJIAYvDTozLBqzwCMgSL+UN3gHompMDwaN/8b6knHoiNwNxsHXb3pAE8GJat+PKDXTPdy7OhIg2q3BB8+N9G/v1QbJZ+nASnpTbEtLSojxPQak9VbxbTwQgGOf9+0v947h2I/Qvu48HekOvInCyAVE7z9aL/g07YsEWujBVSfM1QPA3h/Sz5j/Hddo+9r8/FlaB00Ny1XNxeWS168vePz1Mz775Cu++uwx3z5+zcnzU7QCrRoK1zBWuNe0jBHGwMwI+9ZwaA13ioLjccn+qGSvKNkfl9zNcw5Lw64Vxp1wFrqDyOIhXC58BwwIMdJ0JLdBPg0gFsKWsagBZwN9OFbAlXOc1Q1nVcPpasN13XK5qrhc1VzWjpPGceZqrh0sVFiJsqpq6uWaZy/PeGK/wZYZ+4d7PHzvAR989C7vfvg2b3/wkAdvHbG3N2UyKn3qmjEByPlgrD6AMQHJHa22ff/6Set4IcqSXkYZTLoXSVjyShWCrzyATtLSf+oV1W3MHvlZg1GxtZyRKH2PRXpAMljc1MgXPgFQwnJNNxodOEjgaRwGAU+zrj/xMX1XuFHDtehB8H1L2tczeTeYMZaFACZiRkI/Rh2RJSMXxjZY10QZ5frsFD+mpg+alTAnqp4+ie/swVdnT8UhS9oSY860Aw19vYmSCb908LmTSyJsrOUcx8Y1nDYVzxYVL64XXC825I/u8uBwh5HJmeQFO3lJIW2UGsY5LY0x+aABP0L5IR6ATISJOqyncItKhkrGxghfX6/4x1fX/NfTOV9qphfTqVsXZa2SYRrJaVrTa51e4EIvbyTZ3KQ/8S+4YjVuKHKbaz66rHps3LmfO0GeoMnuvRKUd18U0wt7AwRFqjGZWtNwssQyGBy26lCnqIl98u/3KD0FGenL+/HohWvP/B1ojsM3sMyTsZRYbxw736ced4SxTw6Yu5Ebn6ZcpuvfsbdqvRswNioGrHXPJl0gCj17Q+wJhLSuMEM3AjBtTwPo8GHikobZDjMaqOHuPvrlF+mw/xDQdCBGFXXJ68Qrt4F6d2HeVTqLs5cmiRALYxTXrNVB28J6U3F9veH16ysef/2Czz97zNdfP+PFs1ecnlyyuljRLhvs2lG0MG5a9lHuWDjIhLu55biwHI5K7o4L7owK7mQZ49ySZwZrhMwIuVZkotjostLGoyF1HRt2QCl2WpPr8RQ+jYQfgVWgjXhfBxQCJyoURjgwwk4hPCqEZlLSKjTtmKpWFpXjZVXxarHmZN3wumo4qSteuJaLBi4aw9x4z8j1Zs6XV9/w7Vev+PU//pHjh4d8/Nfv8ZMP3+Xttx9w/+4hu3s7lKX4Ne2OJcQfYyBxgc9105SQqVcYYnp+DoI8xrT0fB7BRE+P0QDoqFBNwmuRP5Pvb7Qg+dwFofbAqzsgvQOhSVUdfw7PX0iVIRjiEcse+kgnRoajoAnt3nYGw23Jq4K6/pA3jZtARTqKMS0Ra4Z+qQmyVnuQEVsYOV7iGHeVR29eAEhxjEMFPT/r1mFX/b2eXMPOCJoAjpTuMRj1geb9KCU+Ae1b6ptmfCCiM8STNhBHlqHj8YhpMVNZl3o2X5lmU6GXKzb6Wv5TPubDQ4OUGVmZhSB1aJpWTN1a5+yPvrXi9/YATCYTa0VKEbV+Rd6gtqA2OefLit+eXvH/Xcz1E8lY7s3q/OjOybTMXxtFWDaPVmdXB6204t1Ggmt8kFNURtGlk3iOAGhFcK3gGkNb+6MpXaecIjL1rm6fBZDEZqpf72k7Ao8Ro3QTvg2vXGAYRWiNImqwGpTDwET3rkMnMSNBAviQ4C6L1lS0liMzDsutqYyaoH+A5DlBwhh4wePHLfFqSIAgQli/S+rXMHYaYy78Kp6G8XMSrWO/74KoeuaWALw6M8KE+6SzEjQQr3PRJvLz7Mc03hN+kibFTTMAXIzIlmTJQFLAp90pkp0+GswIoS+e+TuDoRvTOBy+nxEouSAsXJjjGIBlOupQENepDv9U6G+4EmNbIkDqPQja3dE6x3JZcX5+zdOnr3j85BVfff6Ux1885+W3r1lcLKkWa9yqIq9b9pyyh+XAGA4Ly8Oy5N1pyYPS8HCcs1sYxpllkgljAyMUS4tQ+/fGwXZB0HUmTq+4NSpvMaja/h6Tznc/A3E/DokmtvS56ISMG1wDDqwK1ilFwAQdSsoNLrc0Y8sjN2K5O2LlhOu65fV6w9NNw/NNxbebmtd1w2nTclmt2CzXrM4XLF+cc/70Jc8//5Y/PvqMt959yE8+fJf3PnibR28ds7M7ZjTKsZm32i0m4JOo+LaUTrAYnfRgMirIuNzkMN1cS8ht8UPrxygCBRWLE6U1GpCvGwqZxHvWM20vI9Jrqp7eoy+vc36nY3lrNIFf25eub9plXTl6l3dP3b1nUgbfJIMxACpDmUIMDMV0ZBaDKiNANx0ACI9J77pXL8K7OfE83i/NQr89tQlANr6jiw2SwIUa0sZjjI/0P3G5xMN/Fze4HPRIJUqvkL3UdbMPYhyOjtcpdWNoAwAI0THs7k70vbcfVnfv7C3PT842L799Obm4uB59uljk7fUSeXUu4+kYtRmaZQFnK8410rZiVZ29ZTL+ouV7AwBVNUZMLooxAeXXJufCFHxx9ZrfXV7rJ03D9f5kQgtVAAAgAElEQVReNXtw/FzL4v/OsuwzVTkqXfO/5oXZd40R54T1qub8fMF4HQhY+1no2EIAUbLMA4Dx6JLpqPR5wl1wWo/mnWg30T2heUuyXx3zWzXEOACJlk0fReNRaXCxuVCRVemUVA8lolKTzvUV640KLN4ZeefWGJVbsg+IgCPWkLoeu3XMoGxQjNoQsBbWsolEn6Quka6de6JFWtDADqLBAmrpNnXVHtl3Ao4oSGNIZnhjAADx0Lh0oSYKzuHxs31f+9CI1Cbp+zHQw9q3ZbtE2okgIN1Mprun64f6/uOXRlzEUEGAGJGuD/HeuGro6zFbre07ImoH2QeqLeoaFosV3z4/4ZNPv+IP//InXr+64uLkisXJnHa+YtwY9tQxcw2HOB5YwzuTgnd3phyVOceTnKNRzn6m7GaGXMSrJW18Cq4LvyPFixdInp4FFRvI0QYLTFCJa7mG1hEsK/H0EKyrGNPiw8ritjuCMS64l32SrziHGIdoCzbhUW2hjYDYyw5jDIUYCmvZyzIwloacRVPwcaOcNy0Xm5qTdcW38xXfXK143TheVTUXVc31cs3rV9ecPbvk8ecv+OS3X3H/rTt8/NP3efTWfe4c77GzN2U8GjEuymA8K/EQnJjy17v7TZjfnpj8I34iW6KfUTFYhDbVLAnvB74TDVH0cT08CIG4DLil7OnGuF9qVI2yUQMdJZo7CdgbFMXPuToPyqLi7ETsLfJmYGBs1Rjq83B7K6YBME57eSthT4jAf6giQXPfGv4k/VJqxEuSgHw/nkkMgIK4Pm4nGv8eADhcyF4RFaz6uWyNX8rwy5XWGxzBE4TqICYsgsGIVjtZF6GXSSBJmBa/LGB59fKai4s1tQs5NKIcHM94+Padi91Z+cfVev7NeH/8sG2bj661ffDFclXmJ2f67tE+R4XIxmY+SN65aIOItakr8ccp33sJYDweizHGGIkrS5aV5Lwg4w9Xc76sGy7KstXdyfn0ePZfnjx5+n88vXj59fHenV9uNP9rY+TnqFKtW549fc0///ffUxRekaC9YhsU4zAWJpMRR4cHlJk/otIrASAIn8Ae3eYg3aEepAQfA2I8AIgAXPAZDK4zlj2JRALzzUgiPsOUmEAAiiYHn/QYuitptyRVcymgiMKSYQxkuLlndUWd85tL4GMpBDDOEp1R0dr297ugqGPTo8CKP+mSRBwj16m9qM0jAIgr3Y7oTh0+y41Pacu/q+jW/fHq7cWkPv/kxsHHARC82TLC2PhJtP36pYCIxZjtyhvQLIAmEM1ChHivIFVaL7A09dwpaENbt1xdXPPkyUv+9KfHPP7iMRkZUzImrTJrlGNRHmSGR5MRH4ws749yHs5K3t6dMi0suVGg9YEDLcGyj8BDPfFYvy9/55Z3FnVC00DjWiqn1M5RtQ1rB5U6anHUTqidj8dwIjSqqOvBkgJZUH0ZkBshFw8vrGkpRChFKQ0UIuQmJ7OQZYKY0J7oHnVBADvFL0XUYIRMDHuZYS+3vJPlQMmqdrxejHl6sebFpuGbTcWTdcPjTc2TynF1uWF53XD+zQmf/eZzPv/NV9x9dIeju3vsH+6xszNjZzoJywIhvEtCP7v/YmCrnzcZyF0N1BLkB/Hsg5bEFMfEMIoAAERcANdtAgA83UDT0ah/RcYQKPhrTmtUHQkE6Jp0GwTueSgq7ITvIt8nxzqbsNSQKtLUItYYvqeG3gMWv9HubR6PSL8vhPTtTXmxB+49Y26zqFfmQQLFfQIk3mewzg6vdWzb0JoAABCMRg9dG8IyBHE29KjfMeWmMRHHacu3Ij5rAumBvwR9YTCcnl7xhz9+zap2tApilMmk1CI3p8+ffv1fvvni0/9rd3f/0XQn/99Xbvyfrmp397Plwv7h/IIPdndYmozGhOBCIxgRgex2S+cvWH7YVsDWhCQSRY1hbTJOnPB4teFCBNndqWUyfvL42eP/c766+h+Fc7UqtfqwYdHGsWpqPv/8Cd88/hZreoLvdx/zJaI6jCKZUNiMuDdVXGnRxAXpVSJ0aC0o0t7dlQHSRX/SvdmhRmmIATd9oFy/30x0J/cEHJMTvEjuIPANKz9aoQo401sL4QR1j6sleBi0d2ulZcAu3YdhpG10WA8dgv6ezv7QOHrfpyT1x36EsfnLn5YWFVgUJ99dRHu/Rhwruy0UB8Ar/SJNXAoKVRPA121us90+11lqHhB5t3L0eseU1nawThviG1SR1uGqBlc5qOCgLtlVZd/VHEvLo9zyk3HB+3sz3t+f8N605DgXoIK2gXodLPwAvCQDMrAGtQLGp+PVhN0Bm4YmvLOtKjabNav1hlVds6wc1+sV11XDwrVsaKmjJysIVncbLdOThFXIAVFHpi1TY9nJM3bynJ2yZJyX5EVOOc7JygIpcjIx2NxSGKUwjkxs4K0Qk+BacOEk1MoL27FkvDMreWd3nwrh1brh8XzF52dXfHY156tNxau64cwZrhvD1VeveP30FY1VNDPYsiDLA6CLHrEQr+BoccbRRmUSFLq4YaS3p42ekW/zQGXqwypvJ9+2e9aqBxGtpKA4enrbxAKP3rVeCfbkmIT8dVpQg97qAUAf09KDGom8Rrq8Qec57W38ENejvUXey6YYKtv3wAOA4QAM5G9S93YZZGfcMn7de1WwGt3zOgja89H3bSdHxIXlROO6gEXTAbYeAFiXbqTEQAfFdM7wdW+mxXFWD4VAqBvHat2y3nh+NzhUW6mrVX11dfG6qqrf/9M//bff/Nt/+x/zpi0eLharw8u1mK8urmVclCyMpTGCWB/Mau2PrvuBf8VpgDHCsUFYi3DplMu6pcms7h/tVztv33/5n//zH/94eXmyvvOzn9nSFHlbmdLvIOKFV9NA6wSbuF1vvEdBjfq1WiOs4oYl2rNHL5R7CCDSk1m/iU2/Rh7XnAN48zEGKA3e7TuI/DR9BoBP9yLoqoikk3YPgnwiMOnZWWOUqkQXVKKYScHFzSqHyH9o2vbQY6jx/JuDFRjHWPu4+YFNvpVZEWBK13JVTdSmdgw1xPMJE8f6NamvC05M7xrq6biRRmIadSlEfVQAyfeEOAywW0utQO/uH4xXPyexn4MnUzNoWNvwzTH6OfiQVUOWRRjLfk9MR6bOr4U3UDQwbRx325b3rPDBJOfjnSkf7Y14dzpmXBYU0lLIyucG+hN5Ao9Y1AQLn4xWcho1NLWjdi0X64qz9YaT1Zqz1YrlumLTtDgqMhw5SoEPbFNRbJGxJyOsGH9mfGaxxqsPI2bAS1E2Syu0OJyDpm2p2w1NW9Foyxpl41per1bUqzUboEJwWIzNmWY5O5OCO9OSO+Oc/bxglJVkJseKw2KwkvVUoeplhqtAHJkR7lrhYDfjr2YHXG92+OJ6yWdXSz6dr/lqU/Oqdpw1lmubscks6xpcQIcqYckDz55OwGUGZ62PeUgiP+Maf68UPF16z+GQPgRCnFCkMU+XvXt5oL0ZZB5J90RCr/5aGv+SAgBJZU1npUR5JN3v3n0t2BS1BwAUjRrtPEhpr0zXkQg3/EfPuyYBKJ1nU0kMDO3r6bwOWyg9mvEKaDAtg9GXlihz4j23SQ8ngpMetMUdHp3xS1wmjlsU/N0IpoF7DOY2JlmnuMaDAunGvtvDQw2uCfOhNcnx1ZJlWSE+SOb64uL8i83GfNE6fuGysrhoWl5XNddiqDFJSqJKivN+rPKDAIBfHo2x9h5H1U6pXIsTIc9ts7MzXVxenlwA7WHbZlmRZbah6DeACJHdVmit6Qa9+zoQlnSaUVEruCzrg5JIMzVTguvRfVqE4LZEyXBY9RPZCLRiaINF6YwZEHyKlqMXoNfatwTfJNsD31AiYuIiF30CTu8iG3J4rKNnvIEy9Q2iW3+PgVndd2+gG+3/2M5AuGH1JgFjPso3TEgY3rgF7HCwfQBh+p5uYtM1y9vap7coeB1uptJ9bwLddOOjW7HdXdO3nkzA3QB+xcGNzL5dV6CtkB4VuV4cSCPQgqsV1wTCUhPu8fnGmdZMm4Z9bTkWuJ8bPphN+JvZmI+mBQ8mhr1CmRnFsEG6Y3i9qFXj01mdCm3jtwR2VcXVZsllVXO1WbGoNixdw9I5lo2ydopzBiuWspiwU2bsFhk7RcZIMnJrKG1GLjbsDOe3iI0rBx7sDscGYkYOfp9z53Ba02pL0zYeEDhl45Rlo1w3LZdVzbxu2DSOq/WaVbNivhBeWcNEhJnkTEdjdkYFO2XOdFQieYbNLVY9WBcEnMOoo8BRiDAxwt4kY6ec8fZszIeLmj8tNnw53/B40/CsaTnZOK4rw9IaGpPTGKGVkCqooCbD5CVmVKB5AACSAu6IAPph6Hm1B6qChmDAoHijAt+6rxdytwHMWG8k3BhgG14uSZu6gE5PH1vQgz4fqi8uATFRoIiLqE63no0lApWUB/2QxGj8uPzl+SHhrwELRRqKIKUPOuzQUrfEqDeCdwaGw9AV0r2rAwlhbrvcnzBUg6wCuiEgwpkE2W9VHy0LCcOe9FEtMYZMWwfrBpoNtCY4rxVRNUWWZePxWID28vLqUmRyriZr28yyUOW6cSwEanrPoXMxNefHLT8IAFhHSKv07fLrgRrWAv2O79aaGIVEXdemnGTWiMskBpFkQjYbk+1N0Mx0a++KhqyiHjGKCM4CRUYxnSB5HlB8an2niihBb4nCLJ1yaIWDDGYoOUojwlIMl61y0TrmDpq4fhp7GCxSSavvXnsLEw9hevcrZjd416Im2X1+P4TuQpxyEyNYkxQVogOqZ3bt1vf7+7agwM0mJv8mjfX/d5f7ZRCPZJV0V7yoTEW2hyFmFZBYTX17ujGNinvAy7cLxW5lIG228W761BCSJJ2ou3hLlbG+IfwZjoWY5IpGIJgAAOcBatZAtnHoomJ1cs3q9MpLWgdWNeTt1xy4DQ9cw3u55a9mJR/ujHl3NuLRKOe4MIxNC7r2rn4FH7RnUMlQk+GwzF3L5abhal6xvJpT1Wuuqw2LumLT1Ejr2BmV7Jc5d6c5eVGQZQW5sRSFZVxYprmlzA0FGZkRMmOwMSUq9jEdDDcYFnpeC7ShDshBxIMB19I4aFSpWlg1yqKpWTYNm9rR1DVNvaGuKzZVzXxdc1FfI3lBWWZMipJZMSYrJ+zt7bBfFkwzSyEGIzVC5QMKnc9rz6zjKM/Zz3Pujke8uzfh9WLN14s1n1yu+WxR8W1T87K1XFlY2Zy12OCdETAZ44M7TN86xk29C7bNhNbQ7euOSIjG79YDgzs9jYFRSK9Jck1cT8CqYUxvc1fJFqFLWP+Pss51X/msH9M/01nvASioxQe40iu8zrsWLXvXtw+2lHPk1wBmSfgl9K3nt56TpBNg20o6Api0DZr0OQUdsT06qKF7x+D+OI6+H6nXEWJTeuNG4pwGcNCBD2KVqU4hkXm+rWLEpzkm2VAS4rFkU9O8OGPz+DkxxhDnELxHfzqdAtA0TWtybcSgcWO7WqEG4m7NIgazTR8/UvlBACAmWUQUmIuya4W9PGPc1FRNa5tNVRZFMamqyjjnRFWNnwL1UZRFxuTuAbvvPaIeWxoTMG4gKAkEbQIjtZmB6Yj9B3fJJhOazNLeGlJ6s6gqVmGvrflwnPGTccn9TCi0oRbDmWY8Xld8tVzxojWssgwlowuCCzMZ+bk3hkLInW4RaYyaDyloBrCtQ1owrYPGoa63IFvnAYCEU9UkM5BZ1JrgujJhC2RP9N1+hxLTeYJCTl1w+l3qnw4lDxWgdODBl7AZrCgx2c7EdfLAzEoK1Ie16RZviZoAhIYaudtoJHmv9G8J7+37NwwS2QYAbitjYFsQxfqS9KO0tx3vC8aafvlI47KTFxxGfbR71jjKSuH1FYsnr3hdfcPq9Aqrjsw5xq5m1m64IzXv5/BvRjm/2JnwV7tj3p6V7OUG2hq09RsDiMNzvQW1ODVUtXJZbbiuGl5Ua14u11xer9jM19gM8jJjNCo5yGccZgX3phP2y5xJYSkLi8mEfgekGPns8LvzSwjCC3SudHPdT+lwCSCOli8xgkVAbBfXkqG+H8ZCAUgBUgZrSaibllVdc72puVzWnK+XXLQt103N6arCXW1o9JL9+ZJ70xHHecnBaMQsN0xz6zcfM4EWwvKAFcO+ydgfGz4alfx0L+en05JPr9Z8uljzybLmm6bipFGuTMZCDI3kVGLIZzvsvP2Q0VtH2P0ZzaSgyqGSuLoj3Rp6XH7rAID2g2UwqMbx8LQdFWynGNWFIdbBkHYno3YINmy1qw6nLZrKoE55BfoO2T89H2q45rrcf8I0q/boN6Zd96HS2/MMYBGx3V2p8YG2N5yWRgIwuQGvW7Y5ffCOZLkxtieVrZFXfY8NIvGQqkjbfuOzbm+L5LnemedPk+352rsGopRwXWSxb1NseZoBg/UAQJO5MoqXCddL5r/5lNevX+OaKmyp4efD9BHFzGZlsW7NyNUIzpHZzC+BId1GU2KsGrsVhPUjle8LADxmdLjGKjEuNcenI90dl3w9b2SxWuYXZ2f794/vP3j87PFj57yjXbFewlpFSsv0aJfjD95iM7XUHZMN0ZcBMEKbZ8jOmLsfvEO+v0dTZDQBBKZ5osOm9n9mreOwXfOz3RG/2p3wTmkZaU2lhhfOsne5gMsFmebMc79QIANE6YVinIpIUJ3y6xClT4mxqmTOYesWs6lhVaOrCrfaUC3WVJsNrmlwrcMfH+wVfz7KKCZjstkIxiVmVKJlSZvltJmhNRH4+B8HXepjWqKLLP13eyJThu/vS2ktiasIsQzi0liLrvO9EOmsENu/pwMm0aqI0HirPQlQiEIsWheiw/iE/tANupQriQBg0N9blJcGiBEBVHeN3sAlCLLwXQRUoop1Sq4tedWQzdc0J5ecny04m8+p53OypmLStOw0Ncda8ci2fDy2/Opgyi8Pd3h/VrBrnD8StK694jcC1qJZgUrGpoFN1bJYrTmfz3lyccnJ1ZxzrWitMMlKjqczjnf3Odrd4XA24WBSMLN4WtUWv9lP7QGGCzQcLbzOeRYHJV7QW9goSUPeJiVND+NpEoEc6cgGrWCImTXkOXmZk08Kdk3GQzJolHnrOFutObmac3Y959XVBVdXL7k6a/hWLYd5yeHOLnf3Z+zs5JRlRpkX5GL9IWTa+mPIQ7DdYT7m8O6Mnxzv8fNlzW9OLvj92ZzPlhVPm5rX4j0CV40yf32CfDvh/sEOR2/tUDw8wu2NqUY5m1xwJqMNgHh4IFnI1Yp0Qq9cEB9Y3N9rgsLpI1B8LFKkzy3QnkTBu0HEesTAt4PbYYnKMXCTM0P8rD6DIzbeg+I4n91dWzFVvrMimngUSMYlBtSldLC9RLFdvDDv2xaAi/bj472+CV1tly61N/h2QrzRdliWGVzojTT/VpfI0iDrdKt/Ir3hELy2Bshdi5xfcXI15/S/FbjFOpq8qFOt27ZdLBYA2d7e0UG2bI8Wm01mG8e0yJllBeu27YIyA12pyG3rzH/Z8r09AKvVSrOdslFBm5AmRFMzbWsejkfMrq758uQkr8Xdf/jw4d9JPv5iuTxbzRrEuZZWfay8GKXJoMqFKjdUcTmLmGrXb77gjKHJLZobxoUhG2c0o5wmWH8itkNysUTiVHyqSqaOce1oxhYdgSkdWav+eOIWNqVhOcpZSM4iH+EkLgPEsU/2/ZOeIMQpxmmwfHwUf1457Lqini9x55dUL0/ZvDpnfXLJ5mLB6mLOZrFAYzS3ikfM1mAnOaP9GePjXcqDGaOjQ8o7x9ijQ2Rvl3aSUxcWZ6CVuHGPC2EF0vNt0MMmiQvYZjtNbk4eC5Z9mpIXxjHGLyC9p0agP3ykf4NoVBpDIRWDjWICVl+CZaVbbcEztNkO0vOE0VtZYV5koNTSnnma6L0PXiD18dXQBRd1gxVSiQKuMQKmhaKpccuK+uSK9dff8uoPn3H2L59RfXuKuZizt6k4cg3vSMvPxuIV/8GM96YFIwuFW0PTBOXpvOK3Ga3JqFphtWl5crXm+cUlr+bXzNsN4Dgs4eNiyt2dGfd295iOZmRFjrWClRbrFt76aWr69DrtLSJxdFteaj8GKUXcGgz5XUpG4p4IyazFbVcHcR+RPx3UDZ2nQ0z3/UQM5RjulhOawxHNaofFes3p9ZKz5ZqLas1v52e461P2RyX3dnd4uLfPvcmMUZ6RWYNVCQGTDuoVSM3MFvxkkvHo0T5/uzfmX04X/PPFkk/WDV+7FS+anKuzM67/sGZ1+oqXT77h/s8/ZvbxO9hHd6CYUGWWOkRoR8+WUVCnAdbcMkaBznuQbTtrk6DM+oA0DR6AlAc8P6tTNJ7gEVn8B9mEIXRWtAPwXROhi6Huw5G7b8J89uA7/dYbRtFap6MVuQEAwvzHZ7YyBzRZAuilRXKPF/Lh03bMV7KwGNNVI8iV2E5JQsLiQVFpYvg24k1lBDfuc/F9Hcl7uVI6sEtDnfe84LdWF1oVbevWXV01djqd7u1Mdj+wrnqvPa+KcdtyXBQcZpbrugpGjEVFVRH3PxUAEBHnnGu9PSG0ztFs1pjNivuzMcdnBcVimdWL9b3J4cF/Go0WX8HutwY5ECi9TFAf2W+gtdBYqE0aVS793CO0RqiNP3hlZYTcGtrMUoddymJev2gXotZZoqIeqeY4KoQmA808ZPPu4hanQmMNm8ywMpZlHjYBUi+gvILxObqdO42QxidKJpC3irQN7XJDfTZn8+qU5dPnbB4/wz1/iTu9xF2vYF4hyw1ZU5NJG5hZcGppDTTWMB8VLGYFdlZi9nawD+5SvvUWk3cfMXpwD3Owi05HuMLQGKExlrYDtcLAG+Bki8D7ovT3xlDT3mPukvvwRC6pByB8J2EvAIkekMCOLjKMZ24n/h1IFDY2qJsEJITGmM4MSADFbQAg5tlHjwja0UCQqR4AiCZv6UWYRquo82UZulaHCgxC5sC26n+7hvp6wfzJC+Z//JLrP/yJ1ZdPaF+dM75acLipuY/yfmn55WzG3x6M+clOzp1CmVGF2IAQs2EsjsxH8FfKxXrJy6sFr6/nnDQN67pBMexPdrizO+HdSc5OYZlmGZMsIzcAda/wotB0TZycZBy3zKDtsZT0j+9S+AKJ1dcr9/QzN/9ONZZzAYwQ8IGnBCtg4zwbYJIzHWXs7M642ziuwzLdycU1i7ri8fk5r+dz7tiSewf7HM3GzMYWawty9YGXog22cYzFMDYZo5llL9/j4e6Edy5X/PZyxaebmqcrx2lbM6/WXC6uqS8umJ2dsfPzj5m+/xb2cI+6sLQiNCbSM97BodoBgC5FLLWqYzCf9lQoIQixX3JKZmjb29XtWBY4bHvJ0dc+UM791SGNix0CAF9J7EwfzCdqOp7t43aNX6pMyMfLUIld9dkB4dCgaHZ4kW+DyzxOetymt1fMcVx8XemzYVv27tm+fSZ1Z3R6wzIYWCIpBvlCiO1g+KwfhmT5IBx0NABkRO7Rzhvh95RREEdm/dHXMStCEX9MtojYPC9Gu9n+vh7fuzpf/FKr9tGkbrJDg9wdl+zmGcUyLHvEwE+n2jTND4J7/5ryvQHAcrl00/FuLWH7/NYpdbWhXS04Lkrenk3l3mpjvr5e7V2dX/1dbsfLcm/3G7HFfVfVh85VqAlniIuiVnHG4WwXHO/T82KwjYITRwO0qjTggwLF0JoQ3anSxS31tBmITADxKU/ebeM6Ikd8AJ0L4ML/Fuqw73ncQUuTmiO4UPBpXRqUw6qGs0suvn7G6stvWT15xvrblzQnpxTnF4zmKyZVw6xxzFzLGEdpohoUWrWsUZYY5iLMrWGdZ6wmI5pvXmCOnzB6dJfJO28xef8dZu89Ij/eh2lBk3sGcdGakkTcGrYiZrthHfzu3XdbvwMDdDEyplcQvRowHXAwGncf61gaRMM+B5HhPaLv7YP0jLIIBNO2JFvTJtc1aXMHzELfNbTZp2Gli0R9pG+agKmQHGLi5YdRCfEjinFg1zVcXHH2yWdc/+5PLD79is03z7Bnl+xv1jxoKj4S4RezMb863OWD2YS3Jzk7WYtxK+/yV4uKRa2lxrKoW14tKk6vF5wurjlbzmnXG2aTMe/uTNifzZhNZhxMS44KSybR1d2CVsGD1MeTBEQZJibliJQo3qT8t0qf+3ZL0f7Xm7JN2PouDVLrqolWZLqhcwAVYigyQ5Hn7IrluB2zs5lxPp0yXy64Xi85my94urrmxWbDzmTMwWzK0d6ER5OSMlOsazA+ZQJcw9gWPJqU7I0m3JuW/NW05Ndnc34zr/h0s+Zp23C+XjG/XrG6mrM4O2fv9JKDf/MR+Z0D2umINrNoRrLxV2+F9jtlBqURsqUUE4Dv7QPvp8uDbrMNALQHpZKOqfZbTxvVDpQMeUcSZRSt4ahMe9qPsUU9z5heYScZUK7rrYb3mqA4k3x8jevjwcMk6bWed42mIHxrLLv70rak1+jAyABm6m3k3K/x+9RcpT8rJZVJJGCInrZvjadK+uuETL032UT+6/jOUtVK2zDZ2T16d/fy6n8xVfHX63n17+xyfbxXV/adciz3y5IdETJtMdoGma2KiBNphi6TH6H8kCBAp043KuIwaIvStC3NpmJc5Lw9GfH+ZMTpxVX2/NnLu+bg8H/T0l7VrjarZXvYNmLI0/PFHSq2YyafyuX/6mSMQgxc0s7llKp6HUzwdvE+gl74SLRWAzhAOuw70H8DVZhYUzEYLHctZa3YyxX1t69ZfPIVr37zCesvnyEnZxTXC2Z1w37bcMcp963h3ijj2Cq7xjE2igfkQu2EhYMrZzhtlZe14/VGOavXXF+vWb44ofryG5ZHXzD64F2av/krdn72E7K37zM6mFEVGY31u/M5CHsZbNNMojBjXzq6SiyDiKLj4EsqJpJbiPggzIPKQAAZhvI/LqhocsV0z/ac2684S/9GYbAW12rKZLeUeNnQHwXbsKQAACAASURBVF5D9BBJZ/OntyZmTHjUx3HkjcNcrahfnLH47Gte/Jd/YvOnr7GvL5muNszWG95za34+svzD3pR/ONjjo4MZBYppN1BtfCOMxUfEGZa18nqx4tvra764XHK+WKGi7E9GfLC/x1uzGfd3p8xGhfeouzYsG6Tb/LZbit90/eyAAP243i5C5PYvkvVO/+z2Pduu2DeUJNuje91AYnPLhcDj2vpddVyFiCE3lgdlwYNyhrZTFpuK5/Nrnl2v+Wq54enZBebimrvzHS73ZjyYjTgqLZMs96lLTQutB00zm/PhpODD8S5vjQveOV9w72LFf1+u+aq1nLewXG+4PL1g+eIEdzFn/G9+Qv7OQ8z+lI0YGmu7zWlUhtq9/1MwAebTWdNxztJw2H6u4ra3nSzrsgaGg+jCaarQi6c+MG1QQ6h3OORBjdO7uqWbKx3Mv3bfbefea1ju6Q65SupI532w7B7+iM92uyQOonn7MbyxvIkHPST4VAh7cETA0Q2D9M6AOA7dZ+3pUZJBIQFKSVtukm0iRcP2s73cCg+p4epiycnk8mB3kv+9W8nbujHvynJ9fzRfje9b+OnuDvfyjMa1SNN0ekxFVa2pnbMNP3L5IUGAjRqWxufjaCtKrUrTOJpqyZEIP52M5HK5pFqu7NnmdHdh8t0FOUvNRG3pkaEmwgo///2Z1DLcA0KiKlCkWzuOeDY2K9b1JoGk9L6ruBd4agcPFUJk2LT4gBmPPq22jDY15mTJ4rMnvP7177j45z8i374mW1TsrCvuVhve1pb3yoL3ZiPe3Z3xcDbmTpExy5SyEDLr4UvTEHKmHafrmueLNc/mS56uNjyrVjzftDxfGk6vVqxOLnn67CU7z19y9Pc/Z+ev3ic72qMaCetMcCZ1QybMnICqodrs+/5dJcqurrak2ugyj65Ek9yP3Fxt9vVoZ92k14ebE8U56YOvNLz7JsCJFo3GJcUw5XpDf0XAl6ZUmk5S+IOfCucYbVrM+ZzlF084+80nnP7338OTZ+RXfq3/fl3zLg1/t5PzH+8d8IuDPR6WFtwG1hW4BrUGbIkzGUtnWM5XPDu/4IuTU54trqiKnP1ih7f3j/jgzgHv7U/IqBEaH8DX1EF5RSUR9wfoZuWWksxpohDCoBKPQvHFbT335o9dvUMEuHWvJkyUlBuegu+gudQrMAjDacBkiM2Y7ZR8uDflA0Y8urjm0xeveHJ+xvOzV5y8+Jb39vb56OiQ+4d7lNOCaab49MEW6g3SNmBLPjoYcbQz4eHOguNnr/j19YbP1zVPm4yLuqFeVTw9vWTy7CV3/uGX7P70PbKjHTYTQyXQJDC6o1/xfChoH5SegnJJHkh/azpTN+cijZDpXNAiIKZLyev4Mka3BiMnnSqJz/WT0731hqLz0U1b14eh19GCHgYf3yxRccpgGG6ggwF5dfSb9KN/b0wbDwaleMSfAp8kAMBfShW39NUP3+ER05v60RO49FmMKbiL+kmFi5Nz8/V8tXs4KX7aXi9+apeVGVcb85aI/M14xF/vzDjMDK8WK6qw7KdisTZv8jxbZ1m+4QYx/GXLD/EAVCJyKUbXzqirtWXVtqydsquOfYWPi5zscJ+d6wVfVY4XTnmF8y58DdOjpt8sxRkigE7XjvwcREEWcudDwMVwp6j+CN4beblxnjpXYwgO1JsjGm+LBOrnNAq8sEt4C2XrKDYV+uKUs3/+jIv/8QmLT74ke33JaLHiuGl4R5WfjQv+blbwizsHPkCyMH5fdBRDG5YYgnQrDC7HxwJMLPVeybqe8nq95vOrK/54NecPy4Y/VTXPL5dcuNcsVzX16SXL12cc//JjsrfukO+Mcfh4Aj+W/Zp976aPHe2+6cbYl9vJXjVhurSKFGBANwfJ9iWDMY6vcGq+C66F5/0OeDH/2ltb/Q5qrlv/j+/1foZUsGjI7e2OQ8aFJaPopg10E/pnWkfeQLHeIM/PuPz9l5z/+g8s/vAl9tUZ2XzJnariA634RQl/v7/Lvz+acX+aMTU1VGuvZAQ0y2lNxsZZrhYVn15c8+TsjKv1kszAOzsHPDra5eH+HjvjEWUm2HYJrg40G63+lK574TOMuP5zsUIBlmn4W+npr4NsMU3QK5VuMrros/h6k3zgJrrr2mKHpLVdtklnUOJe++l94oGQepe+P3im5u2pcPedO1wczXhxecU3p1e8qGtePj/h8HzBw6Ndfrq3z3SU+02PTIibaNfQbti1Ob/aNzwa3eGjswX/7+sz/kdV8flGeK2W2p2zXvyOF+fXbE7POf75x4zevocZF2wy8WnMNwBOWPdPUkmJyqK/g6jWB4cQbQ1ar7j7610yUAIENSi8yD8S5GlcBlM3ZNf4t4tVpPOQAky9bRKjNAh/JxbBoJotb2R/jO5tz9KNx7C2gZa9UReabm5u+uZ/R4mbWQ3pWpA3SKVBH6LCCs8OTzmMPOQDxLNWyZuVKVdrKaq17DvlXm75eDLh57sz7huvj9ZVzXxThTMEhFFZrnZ3JlfTab7gfxIAoECT53IlxiwcUm9aVyzqhmWrqDGMnOOuQDEeMS1HPKhVvmyEz9YN9bJhhUYjEcFgXHfm3IC4u9Sx8KcHcV6wpEFngyIJsRCBRJrfGr/rGbPLQY9KYLvC8JwQ9j1vW/LlBn1xyot//B1X//RH6i+ekr8+Z39VcU9b3i8Lfjou+dudMb/cm3B/UjIyCtrSuoa2baibBm1rXMjPNmIQYzBZjjUZuRVmmWVvNOXuTsn7R3t8eLXi16drfr+s+PJyzouqZr7acL5Y0KwXHLZ/Q/7uA9gZsxGhkZ5hPOpNlEiHVrcskEG/byeAG3JCtu/wzPJdVoDG19xC1vGwlduAwwBAbDXVV9fPYbqU57/XLuJYknf3KX6QOSWvlex6TfPsFa/+6fcsfvsp1edPkVcX7C1X3KlrPsqFf7c75d8fTfnZ3ogjqxTSYFrvlldrcM5SO+FiXvP84oxvLi54UVc0jWNvPObdwz0+3NtjNrKMM0OOC2vVwcvVLXe1yUAP+eMmKNgqqfUzyP8Kod/dIA1Msn7gZPtiOtrxntug9HeU2941qDcKfGCwO1tirrnWZ52KgDhKaygzw3h3zN5kxP2DO3y1WPLs5ILz1YLLF0vmJ5e8fXzI3b0pO2VOZtWvt7qGrGnIrKWY5ExGh+yVGQenc3bmNX9arXhVN8xXFXXdcrZY0ZxecvwffsXorftkexPWhQ/g1UHEeiwm6Z23PNIc8jhmf05hbY9ven+0VY0mcN70QCE2yITP6asV7131RlEiH7SvN4Lj/u3JXwMelG6K0nq26xhay2l5A611gkcGd0Xyiyrfv+77jWTnxVC28cebPvSgKbRnmwuH9/q9QGZquIvIW4LcKXLulyVvjwreKSyPMqHUlgtVruuai6qiCcFnTt21zcxFWZarmw35y5Yf4gFoxuPx3GbZRU2zqZ1OFo2Ty8axKTJGAlPXUgqM85xZkTMlo5EVr1fXnDrHJkTDxGjXjnjpSdsPcroxRQz00gFFx93pB6m5CXmYRGP5CFohbuaRysOI7lxCoRo5JaDLzCn5usG9POfqN59z/l9/R/PZt5SnVxyv17wnykfjgo+nE96flHwwKTkuS6xYLtYbLldLrjYrrjdrqqqmaWqc85tjGBHyLKMoCqZlyd6o5HBcslvk3JmM2BkXHI9G3M+WvH2x4L9dbfjtasU3rxpPOCiSFRwZy+i9++gsD1HmUSF3NkL4fyufmb7f/ZBvxREI3bPdSG/VIdEfFtzuMbUzFVo9kB+KsH7+dMjEcvOeqLDjJwlriG/uUQoKI9ikowuLYB0UlcNeLqm/ec7JP/2Oi3/+A+3XLyjP5uytNjxqK36RG/7hYMKvjmZ8uBcO66k30IaUL7G0JuOycry4WvLtxRUvr65YrjfsjEvuH+xzf2/Knf0Jd8elN8tc7ZV/E6yHriOpkE0toNs25/kOwddJ5W1pnF677bn4TkkUtwQtov3zA/zxpvq2r8ubn4mEovY7+hfe7QBtwRpym7Fb5sxGJePRiLtZzovznFeLK15cz7l2LS9Xa+7v7nF/f8pOZrFGEVeBa8lR7uYFvzqcsZPl3MkXHJ0v+e1mxfPWceFgXbVcLNbocsPdv/855YdvYY522YwKaiPhMKDUQBmCM1FQJwPL3ReX3H9zLm9c2brQ6VwNe0lp/7mLxRDYXjrzoMTDgO26utdo/23qi6LjuyEs6I4sjuA6bU8ApdubAqW1pN+YUM9tnY2brQ319zbS0JsYNUrDLcXvRz7pS1T46ZMd6E3mOCzDeFQgARwohWs5EMP7ZckvZgWPaLmb5xznlgMcE9fSqGOtjvO24UobyEvKotDNen22Xubnk8lkzQ0G+cuWHxQEmGXZwoh5jph5I2b/yjl5uWl4WJZMgbG2jNuWslVMYdC84HWW8alC3rRI2Z/D5zMeTBcEdrsIkxT8bZXexS3ppWR+ejeZjz2IO9KRgI/QGrr1463hjspBT665/sNXvPrPv6b+/deMzufcrRo+ssIvZ/8/ee/1HcmRpXn+zMxlCAR0IgXJZFFnFUt3VU2L6pneM2L/2909c+ZldvdhprtEkyxqJkVmMjWQAAKhI1yY2AcX4RFAJskqspp7xs4BEIjwcDc3N7v3u9fu/W7M670WV0KfngCZpRymCdoqThYzjuYTjpMZgzQjyTXGVN6J4q8vJZGn2IgC9lsRz7XbPN9ps9uOaccB10KPvb0uz7VDtoIp0dkEkpQ7ZzD77D4DJJ6U7IQ+0Qt7OCnRouQPE6sLFIrJLeXS7XhRKeZzIKFhINShhMu9ANZh8UUiuzhvc4yXSnkJGMTq9Vf/FH2vT+hWvlOfuA66Op9C2OyxZwW+U/i5RfRnpHfuM3jrA07/8B7y0QmtacJupnkew0/aPv+01eFnpcs/FBqyvFDiJdlNZmC4yLg1mPBFf8DZIiH2FC/s7PKDzQ2uddt0IgEig3xW7u3bpTlzUaut/4uUw9eVDZWyrgazEQezIjAFNWkP5fit7aMW5ZDLflP1e12Jr/fVcb7va4ut+rc+3Zo7dt0720xJtIX3RKBRSrPn+extt3muHfJk0uXOcMq9yZjD4zMeTRNezra4vhGzHSsCFYDTBSmTmbLjhWxsRlwOfQ48j05/zCdpzp0F9I1jvsjonw6Qkznbi4T4xovE+9sQBVhZANjl9K4UbOM2Gt2uGQBX1N8F6+7rIgCW00hA4xHZUvlWsrZMxaOKkam27sRSgV9wadkYd7GyBUdptJXGVeVpqztSwvqLQ/VX7qsi6BKsjtX6dGnKhXr0zp17NVugrvDYBCXnjmv4oys9Un2/Sn2mAjENLgJE3QHhLL61bCl4KfL5Ra/NNZ3StpbQ5vhlOnCifAbGcGw0UwEq8tna6rrFdProST49fvTIz581Wt9G+yYAwCVJMveV/MJ58sSG4dVBknJnnnC126YrJB0EvrX4zpKLnA18OlYTO4NXuneRlqrIxZJb3pXyqYGqyj/PyjQ6NyuaE6Sxpoo56WpEsCxduby+Kyk7a0pvSpYnU0T7j7+4z/Ef3mfx8S2i/pjLSc7LvuKnG21+tttj2xNIaxhnOY9mM/qjIdN5zkTPSVyKkZbA82n7HnHg4YkCreQuRztL5lJO53NOJ4b7SO61Nnh1d4fnd7bZ6rRoBx4vbLbxgpBASdyTPjpZcO/MkXxyhzMhEXHApV6bcLuD8FRBssRyXEW5h/6dQspnNMG6PGxYR2tg5emtKREuvAKlufPU+xTOlTEdjjg3uP6E0c3b9N/5gNHb7yMfndCZJ1xOM16Vjp92I/7xyi5/02vT9TTYirff4bwQLRTzVHM8nnHr5JTbgz4psNfZ5NXtfV67tE038PDQoOcFC6BrpL9dOMndBf9eIAEvOnblozWlUkVgV8pHrn9Jrv2sm0qOJeOgA9mIQWjqsTpXbg2RV1ZpbX2yBBnnUj6/aj7YlT8FCVIKIgel6LRCWp1dLu3ts33U54vTE05mI969O2TY6/Hq3i77m22i0C/SLI2GfIGvNM+1IjavbtONQvZPzujMcr5ILI+1ZpJlnPzxI9IkYy/L6P30dVqXtnFByc2BKFg7VxTeefB2Xt0/U9ida+eAu6AmfKpc/tIVmVCqsm5EpWYdSy+PK7OIzpMFnefda4C/C/viIVbWsWM11fPCO6lfmRp1CJR99vOvPCnVDFuWWC6I2YSwOFtRJVcbjEWrywmLqu9LRFHPaLHsXT1Fm11ekaUN48WBtJZIGXoYdqxlL88JrKYKVVxIj6nweJxkPMktU6Eg8N3B5d1kthjdOj589Pju3S++N1kAANy/f39x6dLzN+P21n2jxWuni6z96XwhLs1Tuq2QjvTwKdxposyj9l0Z/Fbm5he2h8WKsib2M4R+JSuaLt9V62LpMBac1x/LB9YAGizTPETj+rI6SXU+B54Ff5Ex//I+oz99SHLzFsEk4SAz3PAlP+m1uLHVZtuHPNc8SVMOJ3MOxyOmiyktYNf3eMGP2I8C9roBO2FIx1OEqoiAyGzOzGhGueF4lnA0SzjNcr7IUh4enXB1nnNjd4sfbveIW4JLkeA3lzooadBPBnhZwr2JYHbnIZONmPZOj82fvoFoezhfoWXz/gvPx78lAFj3oC1b1asK/3+VMFx/2M2HV/5ykibtR+HBLnL7Q22JFxkcDxm88wn9tz5gcfse/pMhnemC53XOj3zH3262+fXeJq9stmm5rEzt0yAlTvkkzud4mnKrP+D2WZ9JNmc/iLje2+T5nW12N9qEUqN0slScVWe+Tmsq/nVjW6z9XQdHlXuydlHKIiVRynqbpipv6pBYWyiConR18aGris4IV4hP4RBCIYVFSIOUxdqWUBS7stV1KQMYbeOhm/M6vQYEjYcEJbBYubkLBmB9MCqJbMEUMRRCZMQq5MZBl0sdn4f9FndOz/h8NuFwkfPKfIcX97fYacWEfoaoKJpdQksG/Gq3xXYI26dj2oMFMst5RIvZcMbsw9uYJGExX7D7qzeJDjbRMiaVDrviMK+UrzjnEShv9oL3vkkrrWZXFKGSzuIZi9AGaQzKOIQRywyolXz3wkoontQq4KuscFEfXP4W5xV6FT2/enS1FC1L1Vz+rh/X6nh41dlctcW71MIrR666EgGqytwl8Cn66ayoUyaFE0WJZVdulQiBkAIrQUkfZFGDxUiJkSWgKGVVkVFcBSkWnZGumbXmaBaxq0ZCOYFyBe+LoMhuTaTHSAU8No5Px3MeZZqp5znPl+n+wc6D+dz/4MmTe4d8NXL6i9s3AgBAbq29GwTq0zw3b849+eJhptUnownbUtGNAqTnaBuNLoWOFOBV6R9lRL4rZHPRniEHV9SAK4R3Ff25bitc+GXXSPsTleeh5BRwRQEPWQKCpmISAnwHQaahP2J08w6Tz77EOxmyNU+4LuAnG21ubLTYDRSZ1hxO53w+HHE0n5HqnA0pudru8Mb2Jj/otNmNJLGvCSmrJ0rAWawtahtkTnLdCM5yx+N5zp3TAUfTKQ/GQ9JkRjqdcOPqAb1WyH4c8NP9LRZC4Z6ckmcp9wdjktsPGLz9IZuXLxNc9jHKbwj5p9tUF8cEfHX7Jt8TT/2n2b4m86VY/7eK61/epWsIjvqFLYpDhdoRzlPM41OevPUhk9+/R3LnId5gzNZ8wTWt+Xms+IfdDX6+1ea5tk/HpWAyXJnXb6RPaiR3+0O+ODvl8XSKRnC5u83Pdre51I5pB5KQrKTorSzeiy2o1ebOv7woGtsJlqWRy2OlrJW+EwLrimqCBokVRc1OKyRGWzKtSa0lNYbcGBJtSLUhM67Qn3q1zLIonQKBgsBzBB7EvkfkecRK4guJkgolVLG2pEZikNIUBoA1iKo2gbOFtVoVK2oGCFagdX1+NdnaKjTp1md2pdxcWRrAoGxOLH32Oz6daI+tXo+bp2ccjYZ82n/CIJlyfXub6zs9Yi9AuRxhDcqkdKTj5W6AH2wR+wp1eIaXJRzhGBrNQufoLGORpFz59U8Iru1DN8J5yye9ZL2j1n3Ldn4xPBWgu/VPK8Y8i+cK5kpPa+QiQczn6PGMfDonTTKEqRR/uUkhYAk8RAn8CvC37FnhPSjKBtvaSbMKzxuqvolTS7BTGFZrx4jmE1sDrWs3X8UN1FerqzJSy/Iiy8IWhF5iCVzAFQScosgAw1YGaLFupJJ4nocMfLwoxm+1EJ0WJvLRgU+mQEswYm1+NadanWW21tYEnkZgpCSRirEKOXQeH42n3JrNOXUOOrFrbcST0aj/lrXmC+fc6PxofPvtmwIAo3VwYnX2Pkr8SLWjg6FZtG8tUnr+XERSgh+yJ8tsZqlAyDqwr55BF6R1PL01jqvH+uuNS+3mr7V7hTfrXaYmhQrVVoR0Dt8YglnC5M4Dpp/fwT08pjdNuGY0N7ptXuvEXAo8tHE8TjI+HQx4NJ1ijOZS6PPjXo83tjd5fqPDbuTREmWE94oysAWlsBREQtENfDZbHrst2AsC7p+F3B8M6M+mvJOnpFLy44N9djbaHMQRv9wWLNKUwcmU8SLh+PiM6WdfMnj1S7pxhB8F5HI1bWV9SL9f7as7diHoaEhXV0dCNU5ZKl7PWULjCOcJ9vExo3c/pf+7t9C3HhEMJmylC140OT+PPf63/Q1+vNPlcqSI0aB1IXCkIhWKwcLwYDDkzlmfs9mM2Pd5bnOT57e2eb4XE1EGmJkMnGZV6l1g8T5rTFbYXlgVqJTEKlUJaaWKEsJCYh3MMsEod0yNY2YMY62Z5o5ZnhcK37oaBCyMITOG3LgiPMFUq6b0G4mCytuXjkBBqCSx5xMrn1gKYk/Q8jw6fkBH+bSlo+1DJ/Do+oJAgVIWYTXSGgRV4aImKKo0hGMlHmFlyZfreSWlde37tUKxpUVvCDwIopg47BJ4HtuB4t7ZKfdGI07znFGe8dLeFluhTyhFwRdgMjq+z4ttD48OsTG0+nM+1gl3Z5a+caTakaYa33rs/NwSvnQF2j65L8lFBQIKRbayDJuEOWtekIvyklZ8IRWYFA7hLIEW+EkOgyHJwyOSx4fkT07Royk2yRrppK66BNRMnLKcR405Vo2lcIU1XnFQlL15FsvoEgvYNYbCKgC7weB57g6bxGx2yTNSHuNWvBRlxIAVCFmGPTeyyKpxctV4VWmIThYAQEqkp1C+jxdHBLtbxFcPaD13QLizDa0AF1QB1U3SOUocsPRs1J80hsWWSj9XkkQptFCMpM+hk9ycJ/xpPOOhNsxCz3V67WTvYPfRYHD6u8lk9PDu3bvZuQH+Dto3BQAMBndmnrf37sbG/nXZDl4eJ9lrh4kWH0ymOGvJNrq8GgZ40mOmAjJp0CgshoK7XyGcQjbQ59c2JP8sxVUJB9n4C+tWWFOUKOsIUo06HXL23sdktx8Qno3Zz3JeVYI3NztcCX0C5zhJUz4djLk1HiGd5blWxK+2t/jbS9tca4f4ODCLkoksL5VBdaXSbSQAZxAiJ1SSPeWxsx1zLQrYD3zeOxF8NhszeXxEKBRvCp/NbosXYg+7u8XdueZokjCdzJk+POHJ2+8T7G8TbrbxvAgrSrrg73X7JqDwgm9XQkeIVdrCEg9I6witJU4S8geHDN+9Sf9//on85m3CuWYrTXnRan7TUvyXgy1+udtlwwNl0mJvWCkQHql1HE7mfNYfc/O0j7WWK+0ur+9s89J2l17LK6h/dUEGVJNXVW74bwLqK1ajyiyuMy2qt0uXvioY51JjmOaWqTXMtGaeWY7nGU9Sw0ku6OeCk9xymjmG2pACRkiMEOTOop1bCsxabFdK2GFFAYKEc6Vnz+Kh8SjYMWPh6CrBTuix63lseYLtAPYiwUHks+lJuoGi60naUhIrBdIrlVOjSNK6p2RFs1SAvrF+S2Wx6jWoxqw8gTOgU3CWUAa82AvYj/bZCAM+6Pe5N59y+mDGVOe8tr3JQSsgVkFJxGRoYXm5pdi9tsNW4LPVn+DPclgI+laQLjKOE4dLci4JSfulqyw6fuFKVkul9rXCXKruN20fR0UTW71DoWIEgXMEixT78ITpZ18w/OAzZnfvYU9HsEhL+miWJ6wyFZqkbLX+bQKRcqyd4BzAcuejA1b7Xz6j+nwlz2dtAJbnrkBHZRQK29gRKVhgV70EzXVUAUGxlKP1bVYAsGGx160RBwOFgPAUcnuD1otX2fnha3R/+Dr+cwfYjRbWX2aGVfwKxUg0NzCWD8wKgRGCTElmvs/YD1DOMrWWI2P5dJ7w3mjO7TRl5Cv8zbbZ2N446W223z47e/iHjz766JR1BfUdtW8MAAAdhuHDLJv/3in/JRHL/cR6Gw9T7eWjqRgnGWebPbY6XayvOJI+UxmgZY4THkIoQBUkQCV703limQvaMxwHF62pVQ9MJTAuXn2O0k1ezkdlHHKWkD04YvbJF9jjIa3UcCAEb3QirrUCPCEYJSn3h2Pu9E8xWF6KI/7m0i6/vrzHi5EH+byw+Osc7/VKeBVxRNkBLGhXoFNPsxW3eOPyLioMmD0UHE6HvPfokFAE/MjzaYeC652YX2xv8jDtM1ikpIMp85u3mL3xMsGVfcI4Ipei4KtmLVf3awz709tFCP5bbt/oEpXlVwmo4r0ilsMSaE0rybH3Tzj+w3uc/fFDzKf38Kc5u1nGSzbnV62A/3KwxW+vbqPMAqGTYi9ZSpwXMNWWx8MRHz9+wmfDIdpT/GjzgB9fOeDKZouYHLJ5weJXKTOK5/mUVJavMQCV1JEgVPnj4aQkk4oEQWIcizzjZJryeD7n4TzlcKE5TTWnec7YKWYiYEbAjJCZ8FmoCCMLz4GVUMUANMu8LlvBxUnpxXJlloUQAikVvlVgDJ41RDYnnue07IKInBY5Gxj2PMmeJ7nWjni+HXO13MoKg5DQE0TK4mOQNi+AkzMFMKjLDjfoY5/ZVim8pAAAIABJREFUGkKi3nMvrb86cNGA1LSjkNev7tPd6NI9POJ2/5j3H9xlPt7ihwcHXNveoq1CsEX5ZiU1O0HAf37hgE4U4B0OkeOUWwvHqYPFrYecaI3Vmut+SHz9ABMWVrYu95SXXpzGlH3W47/gdfVSumKrMkwN+sEx/X99n/4f3sbdeQSLOUXddFWs+qbYqYMxq9gQLkAmFaAqO1sV5Fn5/GltCRZE/RzKTIMqxRNYZqMUYKQ41iz7U8bLrPbsIgOuAhTFRkax/VdeowwkXPELlADINc7ujMGOJkxP+sweHrFzNmbn7/4G/wdXcZ0Q41EwPJZ8D6uelGZXBLZcmxPp8VhIvjAQa0F/kfLlbMatecq93DHyBN5GbLcPtkadXvzuZ59+8l+fPHl8B1g8Y3C/1fbnAAAePnyYdrtXbu5djv7PVuRvzEh/k/ne/pPEhLNMy0f9MZupIWjljLTl0FkS0UjBKFH5ehRrpQfV+lys2wUusxpEihUP6dPW1cXvFw+1qPkOXmbRZxNOP7uDfTIgnKVsOXgu8nlpq0tHSSZWcG+Rcm8ywzjN81HEbw/2+OnuBpc9C+mstPrL/U5RodlmR5qQtSG4nCstSEfLC3lpq40Ql/nD3cKae28wxo9ifnKwged53Nju8WAy4/F8zniRcjqaM7j9gPil67R3txG+D7LIOqvThGrQVaZk/lko4Nn5y99Oq515X+PYajKUjk1bKP8wN0TTBA77HP6Pdxj964fYLw+JZprd1HCDnH/otfj7vR6/2Oug9ALyIgXXKR8rfaaZ4/3jAbdPThgvZuy3Y17e3OSNS7v0YoVv51B5Cyifd9X/CwO/vsY9V8MqJU54OBGg8UiNR5JZHqWae4sFX84XPJovOE0y+toydIIpHqmMWSiLRqKFIscjFz5a+uTCKwKiKgtZiIK8r64u2GwNF7GVxcCKwhoTQE7hUlXCI3UeU3w8LBKNcprIGVoO4kzT0Yat8ZRdOeNS5HOlFXGtHfB8x+dy7NH2FKHK8ZxFCl2n+NVKfKWVjIErg7WsKLFqfTYsZ6vLW3QEynCt49G9dsC1OOKT4yMezmdMD58wyCQ/2tsnDqIiit6Unh2x4Kc7bYSQtNSIYDjn80TwxEHy8ITRHz/gSyd44T//A/HlTegEJL5YKSJUtYtScKFBdtq03FlS/hbVKgWxBnM44PR37zH8wzu4e4cwy5DCQ/khnh/g+6pQXCvXcrXBsywJTJ0ptGIwCVV4KGvAUjBoLKsaFq4N4arNVVuLt1rMlWDDlQFghcduiYJEXYzHLIVTBQCkWOp416D3riK3ncQJixTFunMl50sVh1Ccriw7XiogVwX4ObBY8jQnzzPM3OIenTHQ70AQsB14BNevoGOPVAickMu+ClvU46rHtPSqCEniBRwj+Wg65ywpquaO0pQzYxgL4RadgKgT292D7WHc8n+fLyb/12ym3zo9PZ1dOCG+o/ZnAQDATiaPh/Fu+E7PQ0Rtf0TL/6Ve5NcH06wzB+8wTYTIc1KLGBpHpvwVwHmxwnCNP6I25OoBLl2iK1t/rB3zlLZSH35lUS1RnAA8ByrVZKdDzu48xE0WtPOcS57kuXbMpShCOTiZZ9yfLRhkczY9wc/2trix3eUglAQmKSz/yoqpLblmL5tWyvpwOHAWYSwSR8ePeWGzw2Rvn8HxgPuzGdtnA17qhrR7PpfjgBvdFp+PJ9zNcvrzhOTuA7KHR3R+8AJeHBb4o+l9+4rxWuvNSjv/3W+q4L7dthJJXKJMYR1KF9H+0STDPjzl8R/+xOhfP0J/eUQ8nLGX5LziDP+01eUf9zd4tRfSERrytDSQfHI8BvOcj5+c8OngjFxbDjY2eXW3xwu9DhuBwnNloF/T5X9BLxuTv2wXgIOysqOTqvzrkUuP3HpMM0F/nvFwOuXRPOVeqrmvcx5pTd8IZtZjLhUL6ZEKDyNVSZm8DPCypQfBogoBWQOmxnw894Sr/1XBiS3Uylo0svjfOocu+eOLrxlEWeVMOfCtIcASO0snt3S1ZXsx49JoxtVQ8mLsca0dci1S7LdC2r6Ppwy+NaUCsktAvbSDl1Z+3d2LTOsGkHSAK8iXpDOEns9O7BNd2SUOPD4/OeN4Nufm8SHZPOeVg1122j6+cghyyBPaXsAPNyOUAE+C6Ceo1HHqDJMHR4yAL33Flb/7Kf6Ll7HdoA7GdbIyWpYAQJz7vT57Sku1fDzCCnwDUWp5/Pk9pp/cxtw/gUmGFIru5gadjR6tVgvf9+sMmOL8S9u36EfpzBbU0fc12KCCeW45xAKKnPplad9q2JdnroqvVY+msYVlZf2yPqEtSnWtxhpQKNlyK2dJz75UEQWIUaUNt7pdUEKLetCqQPSKVrxq1jqSJGE0mjAajslnKeZwwOiDT4l3twl7XYJwk7xx/8vn0ny1BBhaeQyNwyxS+hh8NJnE5b6PC3wT99rp1ecvD4XQ/5oni/+ap5P/cffuJ38113/V/lwAAKCPv/zyJO31fndwcG1unL3rt7xfu1C+YXJzKU11mGdWpdaphfCElucYRQBKwVQRRdTOAWj8reppiyo96YLF3dSt1USsn3H5HVdqv/Vl5kqUWFD+WpgvSE/6ZI+f4CcZHZNzKQy50o5oSUVqLE9mc57M51hneTkM+MVej8uxInR5wQ5XlWut06BorhBqUHBRdHcV3ewcwuYoo9jwWry8t8fnc8tngxEPpxPuD9q80unQUoLrnYjXOy3ePhlxmGqy4zOyx8fY4QR/s4NUzfI338SqXuntmq3/XVn9f34rdnvKPH9tCWcZ9tEpg3du0v+X93D3T4iGM3bTlNcw/HazzT9d3uTVbsCG1JAnOOtA+eROcThN+fRsyAfHxyjjeGlnh1f3t7nWC+kqV7j7TcXZD7WpUrWVIS4neBWU6tbdmRJQuDLF0AiP1AkeJ5ZH85QH44wH05x7Sc5RaulbwUAIRsJnIX2Mp8iFh5aqyMIRovBErAQNlii89qBV71WdfdrckMvjBQVQqVIES8HnXLWSK3e9KI8rLPBE+khg6ixDa/CtJtI53dywmWj2ppor45QXfMmLvRbPdyMuxz77fkCgLJ7TILIiOM81x+wimbm2rmq3beP5OFsXWlLKseFHvLizQdvzuHN6xu3+kD/1DxlZy439ba5uhoRKFVtDNqOnAt7ohSjZwxmHN074PDPoMUweHjL8l7fwQ8W2LwleuITt+OV2nCtLULvScm72VZRbLM21VfTXiuo+QOHwc4s3njP79DbZwyOYJSghafe67F7eZ6O3QRiFJelXGcQmyiyA0h5ZeoDKq5cMjCuKfMV7UDzrp61856psgYZMd44qBmaFKEiUMKNERYW3YAkAKpBErSOq91fd9/XcbCrm+n7qCxVnWZsWrvyV6Ry/FYIUnB31sQtN/uUjFl/cpf38FYKdHokCq5YgZFUWLt+v5lkqQGCdwRH7vg1avtnotnTcbU2COL4fRurddD77f6fj07c++OCDhxRZgn/V9pcAAAA7Go0Go9Ho93t7ew+3t/dvRa3ol/OFfsNJcZnIv2S12E5SF6Nd+bgrZFkMUjOupZaNZXOuIq4pLZjaOmkGtJWuHc6LLlfB7bIASjEhi7iDc6rMOZS1eNpip1PS41M4G+JnGRtWsxfE7EQ+EsdcW07mCZM8Z8vz+GG3w4udgBZ56bpfc/cjWN1TqzrX+Li2YtbftwiT44ucnVaH5ze3OFqknC6m3BqMObi0z2YEu3HAC52I3bMxHW0YTRakx2ekZ0P85/aRTpWOObFkr/wGCrwORK+7dxEQ+zduJcKXQGAgSjTueMDwwy84+d272C8eES4020nGD4ThN12f/3R1ixu9kJZLl89OeRgrOZ0s+PT0jI+HA6bW8outXX58cInLvZhQZEXxn8rLU0etVxP6PNhdmizNz8v5LADlgwwAxdx6nGaOw3nKh9OET6cJt2aGw0xwJj3m+OSeTy6KynSmZCNcErqUtJhCsOpWbQ7W+vNr9GtlIa4dt/J/Yy2KtRd1ypYrZbDCuEIBptKgnM/UBIyd5QTLfWf4bJ6ybTKem2temSS83g55vRNzueWzEwaFAhalt8VWQWZNAPOUtoLLxKqwsGVsgDW0vYDr2206vgIn+f3ZGe+fHaOdQcldrmy3CTxdxAWYlA0ZcKMXI51Cu2PsVLPQKdlckt59zNkf30V1I7ZCRXhtBxcFWClLnoBSwV7Y2fMv6yVnC3klc40ZjDD3H+FGY7AOPwjZvbTHzu4mQStEVNkhTiJFaWVTFlerEX31vMqCOE1TzS0VeT1jnrVd6ERdZ8XR5BGoDL7Gc6jn5PpNFk3WWQqi4Y8QVNsNy67IxmfLU7rqEk+hCi/uqQAsURgg/Q2sscyGMxbTOQxnpI+PSY9OiF+5jgr9FRzUfCRFK+djKYeUUrTakdvuRjoO5UxK12+3w+ONjc69MA7f+/jmh78/fPDg5mQyGfJXyPm/qP2lAKBqycnJyRcnJyf3gH/e2tp6eXf30g83252fJ1r90g6T1xbjvFUF4jhhsLKIyK8qVz1t7ZbPDydkTfTQXMgVG9TFrRSurkCNRS2A8wxnouyJsBbPGBbjCfOTPmKeEueGLeHY9RUd3yczhrNFwiDLMM5x0Ip582CHlgSZ65ohrpY4JYnKOcuwyXpYz9QmO1xjBFwOJsHzI36w3eNwMuXmdMiXiwk/mCXEXkDLh71WwKUooJVrxknO7HTE5PiMncwgQ4UUpRVxofD/vrav2deGK9W3jji3+P0pJx98wfG/vMPio1v4s5zdLOEVcn7TDfmPV7b55W67oOXVSeGOVQorFCejGR8cPeH2eIhSkl/uXebXz11mO/YLl39W1AAontkaaIPGRK0s4gss62ruCg/n+Tg/YGYU08Ryb5LywXDG+8MJnyeaIxR9GTHzIhI/JK8CnS4KLqys/xVzZ22BiYvevwi0ND8rz1d5DcT6d5qtYZnX9d9lfV0nVGHuKENWnkI6x8CG9POMwzThy3TBR2czXgo8frLT4cdbG1zuhHSCgJYyCJMhXF4EarpmxPkFrQ4GvOgzUQK5AswJP2Rvo8UvvZhExHwyfMwX/SOcyUBd5upmgHIe0hrQmpYn+fn+Jjkgj4bkowSbLDgyoD+7y1k7REjYD94kuryNFQohy5lTW7hPH/n1x1CQWTnINIuzAXY0gjQHJEEUsbe/SxipYm+/IuERPkt3eMUFUCnOaioun/ESyzU0nVsWUFtGwq+19S2kxhw5f4/njYjl9m5d6Lc8bbVvX/axCVyAJhBt4rxCv6z2sk7oc3aFdywIPbobHbrdHtk0xWhNOpyyOBmyneaodohTDS6BtQsuARWApdNuu8tX9mfXrm4ddWL1yXjY/+To8aObt29//Onh4eEtYMxf2eW/3r4tAFC1HDgdDAbjMAw/M8a9E7W2Dttx0BtM8xdNoXdFJUyesVyBpcix4vyRwsliUkhRG1XPggEX5a2uegCK/X+ZG/LRlHl/iMotbSvY8UO2fR9PSGbG8ng8Yp4nREpypdXheq+LZxelIFpX9F/jJus7Xb/P5gLJUS7jcuRzLfS5KxVHJuXedMyVVpcw8miFikutkNbpGF/HpJOEtD/BpRmy45Xgx60v8f8ftK+aKUUTzuFZR5Bb1GDO6IPPGf7+Q9LPHhAmmp0s4VW34N9vd/jH/R4/3YwgG4POC8GjPDIrOBtO+P3DI44WM3pRyMs7W9y4ekDsUQQI2ryRV32RJ2RZ82Kth0XKkagUqIcTJamQ9Bllkg+GCz4ZzLk5TrmbGp5YnzMVMVUeifTR0sOqClSo5Xyr5lETONav1fm+iMYxVfRW3dZSRmW1NyvAqbVTPe3ZVNdvpIvVlmYTmCyL/ljhSIWPForE+CysoW8N9zPNzeOUP47P+OFmxBubLV7vRGz6MRGqCBbUZV2GJtA+F1/RCHAUjevXA1JyZmgNwtEJAv7h+h67R5aP+33uTAdM7qT89voV9jptWtIvQIAxkM95s9cuCJDEEHc2RRvJQDmyT+8xkZIo9OgFPybe6ZL6ClTh87VlgLR8hgyDZmBgWezMGNLZDJsV7IVSCALfI/T9guW0tN6r3VeBK7a3rCszPkpmx3rEKg/B12uVcVadQLolHq2npavgTaNIeK3cLzpnyVcqwDi7gm+L2gVLOSnqfYRmCuAyGNwBwtoGvCo8BEKKJVdI5aQqx8iXHq0oZiAkxkI+y8hGU1yaIl3MeXrs4r6lrbgRHFUQ8P5uz17a27w7Hhz9H4NT/d9MOn08GJxODw8PEyDl31j5w7cPABzFnNZHR0eLa9c8I/3olsn9YyXki00fR+HUt+uem4Y4WfO1NL65rCQolmv9K7u2KqjPT7+yulRepIPo/gA/s0QGNmOPDc9DSZji6C+maJux1YrZ7cREnoSFLpnNmidvoNWLRgpYybE9d1zZ51JIC6cJlGU78umFIU/yBY/HcxabMVuhRyfwudZu0Tk+I9aGdDJHj8bYNEO61l+m8p9qiF808t8SuHjKaVbqc1eHOfAtRJnFG86YfH6Xkz+8x+zzuwSDMTtJyos25e+7If+0t8GNXkSbFLIFDgWeT2Icx8MJ7z14yHGS0mu3eXV3h1d2emwEDrJs6XpeEyornV73E1ZNUgqoIv/dioDUSfqp4e58yifDOX+apNxNJYdGcUbExPNJhMQohS0DA897FWCZdVC9LZr/XLycxPphTfDqeKqr94L96dWTNsBspeyf6jYWK38Kz4DCCo/cwcRZ+kZziuYwyXlwuuDzScLtjs+bW21e7IT0Ap9Aekhdjr3Vq31YH4OVtuYBqQGARXmOjSDk9f0tCBQfn/Q5GY/5490HvHn5Cs9t9ugGfhGTkKe0PMdrvQhDj8xoFsOM24nj7GzM4tZ9TiMP0Y7pvPkKbquLlQotlpC86OmyVO05Q3p91JzD6hxnTD3OQhQK30ERNClKt75zOG3J05QsTdGZxjX29WoA0HxONTvjRdJyyTCKqAyw4tm7qugOgKu4JBuxKE0TXTTBQLWuirRZUaQ7rOiEYppWfC6i8YiXk3lldbpiU6zyWgil8KOAIPCRnqqnpnOU4E2iVOndMgKX5tgkBVMRJa+v97Uhqq1RjR8IGwXy5PBe/+2PP/7Tp8CE74HSb7ZvGwA0m7PWJmmaTPLcTIWoWJ6rHf3ivwscN8t/14VVw+IS9ST/Jl1af3Ju7VMBOsdOZzCZIRwEDrpK0ZYSaR2JtSxMhiJlO2yzGweFQjC2zjktTlYiwWdev0KTa8K7dt9WgVyOyl0nMXQjj04rZnG24HS6IM0NwgnayuMgCtjC8ETnTGazAswkCco9ffJ+7ZF76lg3he13Rzi0mjK1VDCF7eYIjMObJORfPubJ795hdvMW6rjPdpLwks35m5bHf7y0wQ97PpsqL9z+woIMSQ0cDqd8dPiEe7MJVzsbvLS7yws7PTZDWaQFal2ZNEVrWB3LoLpnWcQSJz2cVOTSZ6IVX04XfDKa8+F4ziezjAdGMhAeU+WTipBcFgl1BcXvOY3NOc/RSsBfo608QHHe4VR7EJrKe1U51wc2v7cez1Cv2waoPZeCttKpxvhANeetKM6QO0cqFKkLmNmMgc54lGfcTebcmef8dLPNje0W11oeXa+FsroIOnO6vHbVoepHrgmNZn67WB7vTMHJgaUXhbyy00MJwWda82AyQXCCQPLi9iaR55ecESkbHrzRC7Fum6keIOY5XywSzk4GzG7egcAjjCO8117A3+qQB7IsPFNdV5SjsRzn9RTdZsVBp6tMIxrP2DY49IsjnXEks4Rh/4zJaESWZIBaeyxN5d94rFWN4VrJUzNPXgRSnK3G2lF5GJZzi7X50wA8zQ+qlKWmMSWq4xvKodEJV2rzZdcLI3NJfSwQStLpddjY3KDTa6P8ZsBq+dOMzc0tNtNY24ijqeWopKq0uDRJK7lvQRgrpJ3PZuMTIOF7pvzhuwUAAFhrjcXqmlVKrI5B/XzXJ2z9iwbQq0S9XPnuOXRcya1ngINzH4ny4WkNSQJ5jhAQ4GgJSSwEWEtiNRpDIHK2fMdW4C2DiOrelEq9SUnbNLfq+Vu+V+eVNnpWuzNFYzAMwuYEShAEAdpJxlmO1gXKDpVi15dsY4lMjkzmmFkBAALrkKVw+6acNE218/1pFXCyBSGKdQSJRj8+4fSdjxi//RHiaMjmbM5zJuNnMfzvl7f4yW5EV+UlWY8DL8Q4jyeDEZ8+OeGL0Yit9gY39i/x/HaPti9AJ8Xx1jWeW7MfX9HN6oX0QAWkzuMosXw+mPLWYMK705RbueOJCFn4IalUaFEq/iapiRMs99NZU6pNQPCMvrjqe+KCw6tA1VL51AK44RVYsarL/6s17RruUemK61SBgBcBgGorpLp2dcp6jEtZICUZJZe69RlbnxOz4MEo5W6S82ix4BfbHV7uxByEIcoDbFps1TRdhCuA5gIwuZKNQbGudbG2t/2IYLtH5CTJ4TGPplP8I0koFM/vbeJ7fjFP9JyeF/HmdgvtBPm9Y9JFSj61nB0LJn+6yenWFtvtGD8K8FWI9hzmHEX6VzzHSicbd+5QsboZDRZMbhieDnlyeMx0OMZkOfUWkrhgPjfF9HqyimBNtq21i75bKeF11PA0F65jOXeApf5Y+/7KlJSsrLfm3Kw745iOZuhUozyP7ma7ESMgGr/L94zFaYtxDkNJgFUfVYGGxv01+1t40ayRtUvqe9e+cwBQVKH46svUEQElahd1GlPxpisJKpxbG+hvo4ulUBQO0LZA1a5wGXlAJAQ+AqwjMxrjivIqsYKWr8qJWQlnVyyOek41BG0tRxtgx0HJwMKyMEoZnELFnlV6FyRo5cgzgXEChyJxBl3mRvtK0fYkbWEJnUGaHJul6CwjsBasOketfk6ffU+bawJDqmEtxlk6R5Rq3OmA4SdfcPz2B4jHfcJpxr7OuOE7/n67zd9e3iJgCjotU/0CnPDpjxZ8cviEe+MhG62Ynxxc5YW9TVqyCL4s6jesZ3WsC86qo2uHAQivSOtTPjOreDjTvHM64XdPBtzM4JEKOfNCJl6AkYKaNrgpAGnMmQtb9fk6Ras7/28TXa9E4DYC6Wqg0CSEAYShzqxpMlmunpxVq796f228VoS1aKyHi46RGKEwQpEIWEhYEDBLJ5wejXg8WfDr3R6/2u2xE4dEnsSzqiBnss1+UPZ9Pei6iT7WLFGjgYSOH/ODSztkRHx4eJdH4wESRxj6XN5sI5VGmAxMQseDv7uyxdl4zEBnTPOM+cwjsYKTtz9B7W2z1W0R+7ss8LFqGVthG8pkBROdG5fmnnhV67OYO9JVDI+F3MyTnNPjPtPhFJPZxjyp5vLTxn31sCWueIox6+A8D0MTbIrzz7j+jIb1Vr6urZVqbl6w5sS5F2U/mv+LusuL0ZSRUrQ6Lbrd+CkW44rApuYPWL9O48pi7UkJpFBCEIjge6n84a8BAL5Rq1FTI5tC4JwCp8q/8ikr4i9rBcB0xWI3psglp/yRElVy6Vsn0BhsyVktlGwwUpV/jSsnXGkF1TLUlfNYlFsGtjS2KuW/XMxFilM5rUpBaiTMlGCkJZOSyz3HklpN7gxCeCjhKGu+IXDLvN/GHF/B3yvcBOUx35gV8LvxETyNJc2KYrEJSipUbVD9Ef0PP6X/zvuIB0eEScbVfMENr1T+Bz0CkSB0Vtyv8jBOMR7O+eP9Jzyaz+i1W/xo7xIvX+oROrPk828Gj620avms3XttVQmclCADUhlykmg+OJvwL2dTPppq7umQUy9kqnwSVRD3FN8/f8rG3Zd/K3DwlLGv5ttqXu36AaxY8ivep+Z3q7lZWuyiUdZ4BUnaJRh2FU9AaYUJChbB+hwN4f4so/cid5WUZM5njEL7HRbaZ7DQ3D0c8dl4wd8ebPLaZsyeLwmcBKpiOCWgqa9TjV3Dcmx6IutL2xIEpIRK8MZel9hd4t0ncHs2YX73Pv/hhWts9yKCAIROQc+RSvLvrnQZY8j7c0yWcB+P5HGf/lsfgic58H+KPdjGhAojyjLCjUC29ZCzYk0YnLNYdFFjpaSjE64i7am+pRACrDFkWUa2SDE5QGEIKE8iAx8hl6nUzTly7nHUU60Yx3OFxaUogPXKpKiA7FqydnPb7KLr1J6IpnJugNYLv9sAzBUQEcWY2dygF1ndlyzVJPMUayyy3PMX6yyY1dQoA3dV49NC+jzDo++KeAOplHTOyqcf+G/bvnsA4FRpvrOG6J7SBCwJc6rJ3CAdqWghv/Um1qcozcCVYso7rHBoHNpBYizzNMNYgUwKZjGsLZSG06WhUSGZ6pzFvSwXSiGAl1uVogSrDeKV8t5zp0icYu5g4QQZghSYGkdSZqOlCDRVclqJVwUI7Aq4ru6padz9eeP611P86+97zhFoRzDNGH5ym+E7H5F9fp9gPGcvzXhdaP5ua4Nf7G2wGwqkTgowL320lfSnGR8+OOLRdEwnivjBzg4/2NuiJW1J5lSNpL34Nl0VjLRuYZZMfrIg85lZyb1JwvtnE/44THg/hYcuYuh5LGRYRPZLGudq/DQfEvBMr4NYf9OykqZYWvtCCJDl3qwsZ70oU2plseaW1oygYGOzNQ6oPXGlZb003CswUXrCKmVRvS1tKYBLgHzO4lqz4Fbs3+bkLYIhtTDMiEhRzF3OyKQMxykDM+BknvCT7RbPtyNioRAiW6YLLgeTcyq2JuhZt1QL40CREkvB8zs9JjimT064Nx3yL3ctf3P9CvsbIbHyECYHPWUnDPnlpQ20UmRHE7Ik4WgkST6/z8RTxN0OW92f4aRH6osiKLCJ6daf/4rnopHRsMKRUuXPV4AOrBFlWYXiGBV4bOz26PRa+H5DDTTIqYq4fVHk4wuKOUCVROdYV4AVqdAyEaqQXcI1gwtX5Wx1Z5U/qU4LrwyqBkgUVOcX9bi4xlmkjK7jAAAgAElEQVSbTbjKUCi2P2ajKf1HT4op64q6F8aaxsi6ch67+vt1JwUlh0KjxyVAXAFnTXAjRBH+4IS01v2vCwAKwtFqhv65lmUliNZ06XfQpChKGCMcBR635M6QY5FCIUuSiwzJMHOczjLmviNeZEhdMYsZHKYkxBC1MSGacqUpkxtWfoGVqmQcRxGbWtC4ajwyPBIcCydIkaROMsphlGgcitPcMnGSXKqCt1qqZVSraGCwpqu3GurvY6sB44pIQzkINATznOz+MWdvf8z85l3U8ZBeknPdav5+M+I3u21e7Pj4NgGjcSpAW8XxNOOT4yGfDIds+gGvbe3wg50enQDIFyxpfRvzr7J6ESAaAK0ShhWAk7JgEhQhZxl8NJzx3mDGu5OUz3LBoYgYq4hEehjpLZVOZbWwvMzKTUMpeFbFzsqqaE4waRElE6AovVVCKXzPRymH8CRKqqIuuvKQSiBLa2cdZzhXCEyMwxiLMQZjLM5arAatDUYbrLWll8vVlunyXqpxbCiP+v0m6G+qhjWjod6yKDyBRgiMAuMkOZLUKGbTjEE+4TTT/GK3x5vdiEiVpb8NrMTXPG3irwiZ6pjSE2AT2kHES9s9cqN5L5vz0WiAd+TzE7HH870WSgA6xZOCF1oRdrvNIs0ZH6fki5TT4zGJ/5Cz3k02rlwhun4Z0Y1JfMhZpuZVsqOwny7K9Fj/gRUOhoYiXh4j8f2AnUt79LZaeP7SAyKq7chS9jkESqhys8eWkqhUhdV6qAPvGuugfpaq0bulghROrNAIL3vsCq8kBXPrEjaUf6vvNNZGE3wujyteWSfQmUEBg8fHBQAQtTlXn2e5k7KOwFgqercECSvpjk1umfreq4JZTiil1lJ2vj/tOwcAzilRmBXr+cPP+lL1ohmhu/xw+cC/veZEiRiVQniFi8wKS4Zl4QwZlkCCJxQeCu18xlpwvDCMEKjc4tmKXasiLaooP6ljWKSonNdLFFx7RxCsxkIUisYhsU5gKYLDFjZnYYoiL0Z4zI1gkBpSk/JonnGGJJEKG4T4UYQXhDjkqtesKWNX//metWW/RMP151Upf2czjt69yfSjLxGPhnSnGVd1xo8jn9/ub/F6N6ArcshzkBKnQs6mKZ+djni/f4YRitd29nh1d4vNlgQzL4q+rIie9Up0laUllt2rH6kEL0CLgOPE8f7Zgv/neMgHc81959NXMXMZkSuvKNEslrZPcR5HU7h99bgUOce1UhPUXAPKF/heiO9LvNBD+Qov8InDGOmDpyTKUyjloTwPJQVSVZSsyysJwDpX5GUbi9EWYyzaWKyxmMySJTl5psnzHJ1r8ixH6xytDc6a0lvQIA+qKVrF2vRznLPKV267MT5VtHlJKrRQklz6pMZjlCacni44Ti1ur8crmyE9P8QXogzoLMeuuuZKuexnrYcy4NfAThRyY3cDZ1L+++MTPu4PaHkeG17ATicqU0Y1bZFxPfbIdzsczhzTWUaeSAYnE2Yff8nx/vtcbkVEgY9RHkZWzpVlRHs9G0VJFYxAiCqK/wIwU3+xMc4NK8DzPXqbXeKOj5TFwVKAkhVXiCy8RGUaoTa2ILykkGFKShABVW6+pQCIAomUAiFlfV1nbKN35W9BYzdmlYugGc2/cleucVxlU9Z7xRVwLZ9bud1krSQr73dlcC6MEK+KFcHKHHTrM7LYpim2PKqbaR5Rjqd0QkohrbX/6wKAoi3DJ9ber3+79cOpFnrlilpaOt8NiY0rlLavEGFQMMLhyIG51SycoS0FoZKEIsCgGBvJwDpmXkDL8witLZ1vRW8rYmfhBBX3RE1CXFlq5SwXoiy5ii0jqKnlUBnrji4LvUxMyizPETgCz0MoReJgkBoeL3JGKBaeh2nHRN0OXhSTC1mHJJwfvu+P8ndrf5sLVZQpQ9KBrw1qMiP98iHH//oe4mhId5ZxOcu54Tl+u7vB61ttNlVaVvYDpwJmVvH52ZDPTk9IdcYbvQNev3ypUP5uATYrLf3SE3Rew6/2sJZSxTaNUwGZCjmeGt46mfJ/n854b6F5JALOvIiFirDCZ5ni2bzZypxZR2oXDVS1T29BFtsUUnpIT6ICHy/wCOOQVisiboVEcYgf+KhAEXk+TtpC4QsJ6lkeSlcqnaX1WQk958BagcsdOiuAQZZnZGnGbDYlSRIWiwVZmmLSDGtc6SFwZaBsCa7s2n1+IzxaAihR5NRriuJEuVDkOmF6tmA+T/hP+TY/3GmzG8cEyoOKtbPaIqlz3t3XuLap4x+32j4/vHqZ40Tw2ekRd0/79LyAOL5Ky4vKzABNR8FL3ZDfXpKcPHzCLM/I5wmDw1MO/+dbbL1wjWijhe+1i+qNUmEEK65o52Tp0REl9nRY1+h7Y/GsGEmO8vlVQKfwBCnfKy1YgxKWQEkiTyCkRYUeUSskigOMgdl4ynyWoLXG9zy6nZiwFYOANEuZTWckiwwhBZ1ul7jVQkqJ0ZrZZIpO82U/q37JSv67FQdQoc9FfUgTABRfF6WjqzCYZAkEa6zjHE4qHJI0dxiTY/Lq+ssxqVVMfQGxHOs1reSWHywp6ZcqaXm8W56nAGlSuAJVfS/bdw4AhKgq25glGm0sdicspnxfOFGXiHbN2UxFufqUvdhvoVlKmBIE0O0gum2c6JMKwcQYpsawhSBWko6KcDpjnDtOU82MmJ5UeNaBKwPwRNXVin64miBlzuhaLERzbTT3uqv5ZIUo+iIFZ1ozzVMCBZtRQOx7IBQzZznVFMVhPB/TaSM3N5BxhBYSK5e2Zj0jLxjPFaKdbxwQ+Je3yhuzYhOUZCXSgWcc3iJlfucBp//8NnxxH3+UsJ2mvK7g32+2+O2lTToyL1n+HEiPzCk+64+4ORySGM2Pejv85vpV2rEAly0twwsVkGPJqOcKkCBELVCd9LDKJ5M+tyeaf37c5/eDhJs64LHXZSIkiays/nUw0fA2VBZNHfTUACHV1+rPNVI5VCjwwpA4ahPFMXG7RdyKCVshQaiQitIqK1CoLK2spTVVssY1d+ma87GSlBUIUKW1hUBaQMiCVAVJTIxzlk3TRWtNkqQsZjPmsxnpImUxz8kXGTY1WONYFvdqWlxriuIr22pqSw7MZQieRBuPaTqj//iMf8xyfnVpgxe7MSFJYV/X2xRrlM719V3jGk0LWxcpgli6fsx/ePE54lxzdzLgo8EA2e7y8/2tgoXPpghjaSvHv7vU5mzRYdJPmGQJk6kif3DMkz+8x147JLzxAnazhUWuVKyrn0VZ+raI7nBop7Gu8gA1wcAFKKY5pSiMDonDE5ZWAJutgG5ceAQOru5x9YXLbG710Nrw4O5D7t19yHQ0o91u8cprr7F3sIdUgtFwyP1793lw9z5hGPDKay9x+eoVgjBkMZtx9/aXnBwdkyfZusZddq2Msl8q3+I4sSbyl/KocsMLpFX1Z0XMtcMIgTaKJ2cz0mTGYrHA2Spmp/CqVp6G4mwXKf8lSqiiH1zlTamCE51dTXapXjTcF77/zdhq/prtr+AB0CwjjrhwTVfLrJZrVGNXuJ9EifTcyje+vVZt+xjAhAq5vYG3t4O9dUgqUwa5YZRbrjhBWyr2O13u6CmT3HGS/H/svfmTJLeV5/kB4GfcEXnUxSKLty5KPZq+bMd69rf9p3fNum01a92t7lZLoihSPIrFujIrr7g9/AKwP8DdwyMyk9JMkxTNelCWlRkeEXAA/vAuvPd9OReFYSR9fGkRWjcoBa2ClDcQx01zqEjP2qYHcMRXCsFGSi614bwoSMuSnudx3ImIlcIIWGvDZV6wVh6576H6XYLxCIKAUlSQGKIeQnWPP4OAv6ntKD07QmhrebpqjZYwM/BqyuqjL1j89mPUbM04zXnDav5LP+JvjsYchBJVFlgMKI/MKk6nMz46uWCRptzvD/jg3l0O+iFKJ87y1+2z4f3WttZbAkpUlftkyMJIni1T/p+XV/xynvNp6XOqIhZeRI5yim6jANzQfwP+VEcjV8qvcxltDRQpUL7E8wOi2KPbj+kO+nQ7HfwgQPkB0vMQnkApS32ssM0GcXRp67mILR3ULubblqAOQRCVoioEWEUFT1CpFUKgrI+PRxj79PoxZTmiyHI2SU6yTNgsEpJVRp4VmMJgTMUxm2Jdey75G8dzyyCBQgpWQpBLyVpDnuek50uWZcl/uzPmnX5IJ1Aoo6CsMQNaj/b6i91rVlcnQgLlewyjiJ/ev0d6Ap8tZ/zm5DmPgpBhL8CXBmtylCnoBz5/c2fI89xwNk1ZJRsusCx+9TH+QZ/JsEMcvYaJPFJZHSHuCE27PU609b7ZegBq/rGvw25x9S1NcHOF0ieloRsFHI1i+qGHpeC14wFvPzxkfDDGGE1PlshkzaUUDAYDfvDmXY7vHyOkYDHv0BE5djWjE4e8/+gur71+Hz8IyLOCoEyITUqyWFfC9KY90JaitWdA7ui+9V8OgsBFKDR1KQBZHdWVCHIDi3VBnjsvVKn11jiv9pMVsr2TW2NqKwDbK+ZGcth6AtoySlR7Sgrsd1/j709v37oCoBHW2ht3EoCz+ltumcY1DogqAG4nFMTewgz+V5rdfdSlsBS+QI66RMdj1qFHKhWzUjPLNWVpGAD3en2G64JlmjLNMp6vMg77EaHUeEZWwU+VClOn4dXauaXmlltmS8uw2w6tabpiZEshebHOOE0LSgt3lc/9TkTsKbSFZVlymWckykP7HtGwTzQZg+9qkRuxY/d9L9s1G8zW9qFAGQi1JZwnXH3yJdMPP0WfXtFNcx4UGT/pRvx80uPRIMIzmbP+PUkhPC6SnH9/8ZKTZcJxb8C7hxPujzvuc7pwoC9tpJNW1PJ1equuCYWVPlrFXJaKTxYb/vl8zi+uUh7bgAsVs1IBqVQO/pd9BtPqq43p39y6RZ2VBa88hyTX7cd0ewFxJ6TTce7Y0PNdnIOQVTCpkxI7W0bsnHw3TbGvBOw/kbqc9vWlMGJL3wIB0kF1SQvSl3i+JMTHdiM6vZL+oEc2ztisNqyXCevVxoHl5BpTllvraj+tq7rfThqY2Huv0lAsklI4K7mgg0WRFwnJVcrazEjKIT8cxgw95ZQkWz3/fQv6RiWjtYK6RIgMoXzujLq8q4+ZG82r5RW/ev6Cn735kIPId6WMtYYy5UFFp+eFYTnPyDKfxdmU6Uef49+dEI8HRMeHlAEUjfDf3RmSindWUfbX5Gfb6mh02pYSQe3ZsXhYIk/QDRQdzwU/9yJJP/bpRc6VPu4FDGOfMpQMQo9RL2DQdXEjnvZZ9UOGHY848hj1fAY9H9/zMIFg3AuYxRKZO8+nbXAu2g93f2+0FXHRWAWiRci2CiLYEdVCUlhBmRlm8yXL5ZosL91RiRTUdQNs62c7AkNdyXC7XttxtmT93rgM10WcU7ScIqC/twz32/cA6Dp2EvaXr15gCTd4rPaqQdmtsvANyv+d/7WE3AM16tC5M2HVjUgXKbO05DLXJHnJ/UBxHEccRzFXRcEqL/hyseZeJ6YrPAJRIo1pxihpA3du7wdtq7e1Adp7AWf5Z1KylIoLDU9WG87SnED53I8ijgOfUCrmZck0L7kqStLAx4Q+8WRI52CC8b2moJLb+NX/t1j/3w+vwHa80oKyFl8LwsyQPztl/puPST57QpDkjLKc9z3L3447/GTSoadKKFK3mYXHLNd8ejnnd9Mpg6jL+wdj3pr0iWQJ2YbmQLe5o+I6kbVNEeGEvwowKmKae3w02/D3Z0v+cZbxFTFXXkSiQgqhaLsXr5F/m9ntCLP6tRPiXuQTRpEDLxkN6A9iOt0Q3/dQUm0B97BssdLtLh9tLJXtLfeTCrb78HbrumZ8TldvW0kualy2brgTwK8EQejjBwGdXsxg1GOzSVnPN6yWK9bLNck6JU8q1MUGcKjtDWgtoNj7vfN3va8VhYKlcHspLTNWlxvWucEYyY8GPhPPr+IoSoQpd5nR3n7cHUNlTZcFmDWeL3hj3Cc1mixN+LeLU+J+jx8dDZkEvsP9KHKCwONHkz6JlVyml8zygjRXpF+9YP7hJ8THE0ajIbnnY2Q78U80/ze4JcZuA9dayrITkNdLDbezG+t8IykMCoMnNC7ev8RrsEQ0whoUBYoCz2qUi1JA2BJlwaNsfhQKaUukLSrjrURQoKr36wOonVVsHfk0ikn9qi2IEa3v1kLX/WicIC6tIisFs0XK85NzlusMrZ33c5viuUtHbX4ndoBSttctYJtCXi2OfiurrOYg2y6a71/79j0ADgnwT1iA64pBHeQBIKu0kTqV7ptuFtACSimIBl06d4+RByOy6ZpplnOal1ykOe+EPXoePOh1OM9TTtYpXyUpdzY5w0gRyQCpLb4tW4u7FQBix83UvnvremWyaQG5kCylz6lQfJnkPE8SklJzEAfc73UYSIeQdpUXnGxKZhpSTyHigHA8JBr1SeXuPd2eqjlBS7P+Psh92u5LJ62kda7/INfI2ZrL333G+tOvkBcz4k3KPZ3y1+Mh/3Xc4bVYuMAroUH5pEbwdLrkw1fnFNLnR+MJ702GHEQK8sr13xCVaDGHa5J6e01KkD4EMQsd8tF0yd+fTvnFMuNLETP1QjYq2AL77FTEa/XTvG5JsjrqSeDO6z2PIPLpjHoMxyOGoz6dTozyBEJtdQRoqTACEGa7jjftPrud7s0qdV1z3b3nSLJlMrWYZJtp1x23X+3MVdIcMfihhx/26Pd7ZGmfxWLJ9GrO4nxBlhboQrtz2wZbvkWkbQ/NTa1eZwsgyZVHKSQa5aprTxOnYBQ9Phj59MPABURWVv31wd92K+usSl0ACf2wy5ujPuvNHf7vp1/ym9NTBoGkO+kTKd9lmOiCu0HET0ddTlYpX56uuMoFxUXJ6tMnvDocMXz0kNAfY6RPJisBVz3MehWstZS6xOrKErYulsPWIGA7T8h9dz8I2D0Ki6ww+6W1ztPUilFtQMVqhYASKJBWI0Ut0J3CIK1TGByaqfstrEEYg7Stgjot3m5vppZqrrXQblGqME3mQbuEcWkFxlrWSc6Liysul2vS0uFxSFmyrYd+HcBnh8Kui6KdfVsHIN7cQ2t9BdjvhzV1a/tusgDqZ/0nL0WlWWPZRqzgLBthsDsWwX9kWK3/K0ZslEJEMcHRIfHrD9icXLDY5Jxoy/NNxrwb05WCO3HIgzhmsUm40oZPZisOJj3CUCG9gL4RWK0rYtoydYtoEZhD6rN2N8ahch5RCMla+bzC47PM8LvpjMs8xVeCozjkbi8mFIKVkbxMC54lGSupsJ6PGPSQoz4iDtCi0l73BdnOSnw/lFTREMtWCCtrCQqLv9iw+vwrlr/7nPLllE6qua9LfhQG/PXxgHsdwCZAiVWK0gt5eTnni8tL5kXKm90RP7pzyCiQ1bmv3tvttrUM1dl764zRHbxKrOdhVMDGevx6mvD3F0v+OdE8UTFTFbKRAVoouJVOKybU5HVXkd312bsE6UmCKKAz6DA46NOvBX+gkFVhIFt7dfawzC225cEWu49WiG1k9Z672xmUlUADRJNm575nqRRxibt39XYd8+JExJYhW1HHnGwtvnqfAQ0arRCWsOMzDgZ0ehGjYZ+riwXL2Zp8k1MW2jHufZjjvXnttjpor/KI2CqQVnrMvZCvCoG/LBByRU7Ez8YBI0+h8CpDsT4SkmzPUP6IRmA1lBuGfsh7xxOeXi15vpnxZHrFMPB5bdTHsxZhDOgNB4HPz4+6/Ha54SIryEvD6mJO+vGXXL3/mEH4PsHBgNJXjRdgVzWtPaLSrU0FcOMUANEant379lb41su2DcZ0ga41qLCq7yFqv47hVoFdKVvuWKIGcFMVf7u9/ekyst4vmn2XuzMWFetccz5b8/JiTmY9jFAVGmedcrsVRA03bJQgsa1q2K5r0Xxul1eYSh+27aO69rwcf7dCiK+b/p+1fasKgJTSGoRtoie+Zhn2SWC7nPbrP/gfbI2xVdGFAXTgERyOOHj/bV58+oRkXfJqueHLJOVpkvJmr8vQV7ze6TDbpHyWrHiZJHziCWS/g40CkB4dMnxj8DAuFqCRsy2NqD5DsqIKRHQ6di4VaxVwKjw+y0p+O1vz1WaNRXO30+ONXo+h52MQnOWax5uCF6VhHfrYyEccjbGjHtpzgqIOzmrWc2dZ/0z0aXeZ2T5ro1L1lAYvKyhPL3nxr79h8+QFwWzBJNvwttL83Z0D3hzEdGXpLDEB1vO4SAs+nU55sVgwDgN++vAe426IT7GtH3+j7tNeo/bmFljPR3sxM+3x+TTh71/O+adlyWf4XKiQ1PMx1ML/BqVr535Vv81zsUglUZFPtx8zGPUZTHpEvRA/DFBKNmUCGu9NC3e9DuqzrfHX5/ZtpdOVjnBV5Kxx1pT77fL6jXGWt7KSpua6cExUCIVQrqqarCA+hKgzDKhSNS3tYjGm0m1U41HY+gwENa8VeFIhvZDQD4niDov+msVsxWK+dJkDZRWxv48hcO0hbtezbY1hJKUUrAnRKNApYpk7OF0BP+t4DEOFX8/H6JtpQ0i2YELtt0ooLZ4nGcURf/nmQ/IvM04XC2Ll0Y1iDkMfUcWdRApe7wX83b0Jr56dsc415XxN+uyck3/9kM7RASqO8PoRpaI6YBHbZ9JA8mzH0SjQtVBt638NKbqLW3Td6jlXz25fZ2xs9pqFUNEMtcehXpmbeLWFW+TfNcHf6qv93o5B0Bwo19Tj6MAiybTgcp5ycjlnkZSU1uGxNP3amxaj7uvar50Xbt3bx7nVnmsCdltxIdWU23UJv6/tO6sFsOtFuX1R2udB7BH3tzKovbtYIdCeRI76DN55xOmjhxRrzXxT8izP+WSZMOz0OJCCe3FIMugzLUquipTHq4QCyOiho4BDT9AzOaEp8WyFEVDz7IpJVZnt1A62QggyIVkqn1Ph80VW8OEi4fPlisxY7oYB7/V6POzE+EIys/BlsuFxXnAmJVnoIYZdguMx9EJyUWLl/qa+QSj9udoOKdSekPr80jEkTxuYLVk//orlh58gLmd0s5TXTM5PI8V/Ox4y8sEzukr5UxQGPj2/4ovZHJTg/cmYdw6GhBQuB7yx/m+z7trXKnx25WFkyEx7/H5e8IuXM365KPiMgHPl3P5WVLDVu3xi29+NyoaprH7o9mN6wx798YDBsEfUDSvkW9EmUmq4XrHzVG2Tr2+wzsGgnVsUXYP4aIqspMxzTJFjyxKjNbbUTvDr0lmoxiAbAasc6IySWOmAsqTnIT2FDBTC8/D9AC9QDodACYQX0OhBsgp2bbwSW+dvs0iVdJFC4YUK5QcEUUTc6xB2I+bTBckywWTaVcDDsusdZKsc3GKROa+EpJACU4HGfF4aWJUolRLYLu9bxTgQ+DUGvK6eT3u87eixWjLWA7AaTEGgPB5NekznE3579oovlwsGszmjOxN8qcDkKGMZ+oq/Perz7GrGfJ6y3hRk0zXJh5+xfPMN+qM+XuShpFdNVzScA0RVendP2WxN262CrQRVS2hSIZQ2z2WXCQhq/8K2l7YnwVaC2GGLtP2XVSCdcPdse4puVrbrLvcs+jotteqzuW8j9GV1RWCspBCKRV5yvki4XG7IWyBD20nV/d0ENNVWnG/mBdJYUBWctWivepUgaK3zmjV6p2gFtH4/NYHvRAGoSdQ12yxQWwzt6GMt4/ibcvd/XduSdnWaJRW6E+E/vMvgxz9gMd2QLhJOZ5qP1xl3koy449P3Ja/3O8zKkt9PC66K0kU1l4a01+GdbsSx9OlLSWS0C6yxLie71mbdbSsilg7Bb4Xk1MBnWckfVhu+XK5Za83ED3iv3+Pdboex58B/XqYlf1glfKU189BH90LC+8eEhyNMIElNjhAOoes64YuG9/552z4lVFu32m8qK0hPz7j86FN4foq/ThnrnPcCwd9OurzV81BllecrPXIU54uE35+fMc1y3h4O+cnxEUNfQFqyLQzzJwyn+sNKD7yQjfH5YpHzi5MV/3CV8diLufRCUuVXkf5t8KC6sz2PQjvQSIBQ4IUe3UHMwZ2Jc/f3OnihjxBUbnUq7Ii29afdNVHvqbpipsFqTZlrTKbRWUmZpugsQ6cZRZJjs6owUlmCdme0wmg8a/DsNorf8S/nyi2lO5bSUoCnqh9X6dCLI7w4QEUBfujjRR1UFCBCHzxZkd52La6RnBDUsRJWOQs86kb4YUDUiYi6MVfnU9azFfkmdxU7m55u4hFfY30JiRawwecCi9UZalEQkeET866VjAOL9CRCGWfZsy9A944jGg3bgilROiP2FO8fjXiVJXwxW/LJxQWPuh0O+x6elFirCXTB62HMfz+a8Cq74mxTslqnrJ+fc/WbT/AfHBNNeni+AOnc85ZtMJy7dw1aVb00rTiaWk9qjpta3hO7n2dv935v+7ANfHNltFSKQwOLK2oUPguijqa3zQnKjifmlvY1ZuF27evsqurTxgpK66z/2bpguilISlwmTGv/NsF9TSyBuGEsFU++ZYxbaI66XsE2oHH7ndaXq2OQ8j/rEcCNreVSqev63Khv2Zqp2WsepG90NXe0YFW5iwylp1DDHsc/eR/98pzl+SVXacrjdc5kNqcnBzyKA/pRwHvjPlm+4bN1wrTI+bTImCcrpoeHvN6NuOP7DD2fDhBag0fNs50mraWgsJI1ihmSC615skz4YrnhNE3JTckd3+etQYf3R32OQp9SWE4Kw+8Waz5Pc15J2HQC1GGf3qMHiGEPLUAbF+HrlPyW5fK9bLsCQhpLoC12vmLx5DmzP3yBWG3opSl3Tc5Pxh3+4v4YjxR0jrUCjceysHx8csp5smQYdnl7Mub+oOsQAU1d2tdumeaNBNXyDAgH71uoiGfzgn85XfI/LtZ8IaMq2t+dNTbunWv97SkBltofjlCSsBPQn/Q4uDNmfDDEDzzw6gIsdidmaSe8bux8aNAAACAASURBVH9flJYyLyjzlGKTkq03FMsNrFJskmDTlCDP6GYZXQwdAbEQeNLiC0koBbGUhNJlVCshMRVIUGk0mYVNYcisIcP9TrRhoyWF71GEIWkYksURstPF7/cR/S6qG+HFPsr3QEmEFDuZfOx5Zhvj2oIUilhFBEFAGIVcRVfML+ekK+cN2DMdYKdm2y2tUjYK6WJtQPBFscG/XNNRHgE+oYFuCCLwoK4SVwsQU2eJ7CmSzaSqoECTcNDr8NbkgFlWcrac8oeXPvG7b9D3AqSuU1AzfnpnxOfrnM+zKbMsJZeCxR+e0HnvEcHDI6JOwEY6xcVNtXLX10cttUy+LsMrHnd93++mtbX+qgLXt+59u/0nap9C64HVS3rtxi2b/Y+wna/j6Y0fou15aXwTisJKFuuS2bogKQRaemiK5mM7bO/6+cbOnbZ+jz2PSJUu03bE7X9vB6sDSQWBZ0T5ddron7d9VwrAtclb4YqmuOJguxt2+4ida2UnCWjfXfBNDG7PYNMIcgEiVMT3D+n/4E2yk1M2swWnmeHD9YaeJxCyzxudkDuBhIMhSkm+TDac5jlPypLp5YzHm4iH3Q53w4BDT9EXikjU2IAGLSyZFSy15bIsOc1ynm8yXq03pNrgAw/CiPe7Hd4a9bgTeiAsp0XJr5cpv14teI5iHQbYcY/g4V3Cu0Py2MNIV71QVuu9I9Rumz98a2mAN1f5u2k7OebmW0uY5qxfnrL6/Ani1SVhpjnMc96NPN7rxxwHAorE9SMDNkbwfL7io4tLOsAPDie8dTgEClfeV7fz/VtDuElo14eeUmH9iFcp/OPZkv9vtuFLEXLpRyRCYdplb2uTHtgJRNtdCcAgfUHc6zA+HnNwPKbTj/EC6eK56joS1tGKy7FvW0KOu1jjzu91UZCvc5LlnGwxp1gsMes1QW7oFoa+KRliOBCWo8ByHPiMA59e4NP1BaEviZUi9jxCoRxjqBBMrYXCWDJt2GjDptQkumCZZ0yzgsu0ZGYNVzrjcp0zX61J5YrUn1J0Ixh0CEY94kGHII4JwgDlK4SULevwhkAxYZ2iJEAFksG4SxAoOp2Yi9NLVldzdFmXJhYtK/fr6Wv7PAS6Qmi8VCGfldBbpHQERHi8jSYC8Grre1/K3tS9ZVvaW4ApeDQZkJYFyXrBR1fn3FnfJRiFxEq5WJQyxQ9D3hqE/HjhcTZPWBUes4sZi0+/IH7rLuPJiFwqdG09IG6e7t64BC0Dx7TmXslBI2pDpP6IbXxYdZAblRfKtJVOSyUQRYtfiB3e0T72acH8tRQOx2v2peP1J9bGg9gKaSMEhRUsczhbblhmmtw6IKCtamabAm43Wuk33PXaAYFl67SrUmybLIC25lp7WcW1w7nvpfCH70gB2OqMLW0Vx9Os8880kZjttiWN3VoA3+zY7LVXWgjn5vEE/iCi985D0pNXbM6uWK4LXpYlv10lOOIa8GakmHQj3lMenTgmXq55tl6zKguerTSzNOWZ8pgoj4HnESkPKR2kZ2lKMmNYlpp5WTAtNQutKTX0lcf9KOLtXod3ejHDQCGE4Kwo+XiV8O/zNZ8bw2UYUA57hA+O6T+6j+kGFJ5ojqIbsKGaZm+yEqrnQvX5b1wJuO2e7D+DLd+PCpDTJcnnX5F88Qy1TBlmOW+g+flkyA8mAwJbVoA/EVpIzlYZv7+YclGWfDAa8eagzzjwoFhXAYJtDbJlgl5Lz3TX3Lm/x7qU/POrBf80zfikVJypgLVUzvIXgqayiai/255gi24rCDcVSLqDHgd3DhkdDYl7AZ6vGtepU3QreqRmgdtFtNqg8wKd5ZSrhGy2JJsvEKslYZYwzDMGtuRABRwHIfeiDneigHthwF0f+p4i9iS+BE9YpDR40tU8l1YgWwABNQSqxqJtlQhmDYXRZKUlLSxX2vKqMLxMc14mBdPUcplvuMgTpsspm8uAZSckGPSIRiPCQZ+gE4PvYgpEdUSwSyZbYSUU+EoiZYzv+/iBz7mC5WxJkeWuvPa1/P2aKdev6wdUz02AkBR4rJRb80+yjOEqo68gVorXbYGKBMKv8uJMBRZ0YzpvdY86k8JqKHN6kc/DUZ+r8Zh/PT/n47MLuv4RD7o+Eo3QBbJMeKvv8/NRh5frhMs8J0lzsi+fs/74C/r37+JHdyiUqx5ZP5mvc3a0Y953DPSWPLKiLcwERriUvwb+uUXHW8tYbGMMW5b1Njix4iEtru0kfy0FbrDibgoI3ONDolpfa53wLxEkheFqkTNPcrJSYKzYei6qBWiEf1t8fA17a9Z259pW4G/LHcOWydbSynmXbKWgODZS/udVAFpOsXqdtgpA9YHdimD7LqQq6aPluWkHs38Trc10bKWMuMhkSx4pgvsH9H7yDpvzK5bTJXOt+TLNYJ1ihcAMO9yLYw5in67vM/F9jnyfkyRhkRdkecEpOZdIlPQQDpy9ymUtXQS20ZgKzqIvJJNOxGtRhwedDvc6EUNfkWN4kRs+Waf8erHhs7zkLPDJezHBgyN6j+7jH47ZKIeCpqrI7WaO/xOC/dtQAmotulL+qvW2DT3UJUIFtqn2t3n2iuQPTyhfXhCnBQdFxg/7Ph+MOtzv+JC7Qj8oj1VW8mI+58l8RujFvH94yL04wNeFw22vhcKfpJA7fH+rQlZa8NHlkl+cL/htJjlREWsvwMhW3fud8/l9eq7vZxDK4sc+g1Gf8dGYwcGQuBsiPacYiDYzMW3KrPUIiyk0xTpjM1tQLBaY+RK1XNFP1hyYgmNpuBcqHsVdHnS6TMKYYejRDxQDX9ETldCHSlCZ7Tjbf7d8ce5PWdUBkNU0VeWBkGyQLA0si4hFZlmnmtNNzpNkw+N0w4vlmouVIJnPSKdz0uEQbzgkHvbxex1U6LmYgrZy1sIFb8rG+oJA+Yz8AUoZ/FCyuJyzSVJsaapaDrLFJPYC+FoCq3luUpCjMAZOtOajtKDrQT+I6AeCQa4JhEJ4rZoeTdtfqz3a0gVK50wCxTsHEz6bb3g2nfKwG3Lgj+goz2EDFCljv8P7w5CXq5gnFxuu8oLp+ZTVZ0+ZvvEah/cOkL7EVJX23JOyt3jWruf87463fim2P1Rpm7caW7V7vH429ZruegBqtavuStQZA3/C1ruZ47SCAAWNcE1Ly2xTcLVOSSqwH1srX+0iYl9/y2oKWwFjqnu1O9giBlYvdlJvdyu8unUU1V/SCuH/51UA6tYI+0b4t1a0CQu2zcatXANN3QVHo9uF/TaaoIapdMMxAgcNPIiJ3n6N8WxJdnJOnhZcWovJc4rFmlyXfDCER3HIyPMYD3rciSNOlh3O0ozzLGdeFqxLzcoYMm0odR3vbogUdD2foRcw9hWHQcC9TsS9KGLo+3hCkhjDSVHwm2XKh6uET/OSM88j7Ub4dw/ovHGf6O4xOgjQwhXDEJ5EKkVbu77OLG5hXN9U291Hze/6+TeWxnaASGvxS4u/Tjn95AmbL1+ipkt6ec59ofn5aMhbXZ8Orsyslc5KP1tOeXJ5RaIL3hvd4fWDMX0fyLMKyPs2zfG6sLMoUCEJPk+TnL9/ecWvN/BUdJh5AYWqAfCr8rBU0f+ibXbUfVdHAxKCTsDoYMDxvSN6ox5eKBHKtgq00PDXNu4ZxmJLjU4L0sWSzcWc/PISsVzQTzPuYng9kLzfiXkUBzzoBNyPQw6CkEBJJJVFSu7WwlRw1fW+s1ClDbB/JLcDulMfi7gQcuoYna706AqPu4GCyIdBzDwvOUkjnm1ivko2/GGd8TTLeHGeMpstSXozivGI6GBMOOzhD7pI39/qTzsWaMWWBVgp8KVkcjzE8wWekkzPpyTLTaU0VYvYWOot829fAtX9S0HpKRbC56uyJE4yxr7gaBzxqCgZCYOHRCgPFxTYHpvdJaPG1YZbzzwlUiF3hn3eP7zLb86e8uJqylEY8PBwgNQaoUs8mfMgVvz8oMe/zzacljmblWDz7BWzjz7j+Gc/xA8VRZVVYRrhb5vpQX12b1tC6/bd3Yj62qKHa4r/NkWwvWZbJ3ct6moPQC0SJaJKXdxdp1295Fpx9PaKbvlVHXtgnbAtgEVWcpVkrDKNxt+ecBhzy2O+QXbcsDBN7E0jj7ZHJbWxev1rFWh9Q7jNoLlOdN+f9h0pAKaKEK0tib0o1ro1ilUFIsJWcdgWBpI3F2X4DzeBkHU+LM0TLqSAQBFPBnTffcTog1ecv7oiKwqurIuwzmcLitJQDPu83ok5CCLGcUAv7nIv11xtMq6ShHmesygKNtpSCKrzeUPHFww9j3HocxiHTOKQnqeItKXUlvPS8CLN+cNqzW+XCY+N5TwMSDoB6nhE/OYDonuHyE5EXoGvWCURvleV/GwBf+yt99aftZ30txYDwBbmpx6IoObTjoFILIGBIC3Jz66Yf/6E/NUl3TTn2JS8G4f8eDzgwFfOcgJQPkkpeDpb8WqxZNzp8LPX7hNHPuhNde5v9wez23amrMAL0CrkLCn5zdWKX85TXvoD5l5ArlSV525bm73dt2DH8hQGpMCPfEYHQ+4+OGZ8OMRIsFI3XhBRcZbanmhijEuLyQrKdUJ2tSA5PcNcXNBLE+4Iy5uB4gedkHfHfd4b97kf+3Ql7sijKCuo2vqsvDpQqC2eBlynVlQ0W+tObOfT6Ik1jnvtCrdACVpVfVX5jCpkGCqGnQ5vyQGzouST6ZLHiyWfLBIeb1JeXG44ny9YLBaEBxO6dw4IR0O8IMRWgYJtjAQhqqw8cPf1BIPxECUUUkiMuWCzytnWva6Z+G0FmOq+KpvV02RCMrUeX5Wa3y43POz4xL5HlBu6GETsu/m1qwe2+76JHkwJKCI/4Mf37/B0ec7pcsVXUczhZExX+VC444KhF/H2sMMPeyFPVjlXmSC9nJI/fkry/CV+9w2QrkaKC0doKZvVtNtAULdMeO+1O7sWLRpsrLXmEwKErCz86r2dNa15R70kYvc34Nz3N4n562Oqv9coABbn+kehrWRdWmaJc/0XFXBxJfuxVdyMqbttaGbPBWFrQS+qI4ua3m9evHZWQYO93Z73vrLpNrWVUv+RqNQ/X/suagG0qLTJXr2ui1XRxlzbS9uHYeFbCQJk12lFrc3WZ0laQOF7hIcjjv7ih8xfnpALS3E+ZSYMOoNNmvGqMLzVKXh3aHitEzKSioEyDDuSR1EMJqQwlsJU0J7CYG2BL8H3pDvjVE5vLozgXAvOMsPny4RPFiue5yWnUjCNQtJhhH93QPed1+m+dhc57FKoWlMVSC9ABSEEHlo678nteujexvjGW80V7E4cUrXSlbxxAsizEJYWOVtx8uuPKZ6dEi3WHBQ5bwrLXx4ecq/XIZQaCgNCYbyIxxcJT5IEoSQ/6vb5waiLb7KmYlsj1P4o7Qhn2auQJIWPz9f8w+mcL0TITAUUtdu/sS7r6P96mm0CtU2XfuhxeHzA8b1DeuMexhU42Fmeuorb1qK0CG0p1hvWl1OS0wvM+ZTuKuGuzXgvkHww6PCzwx7v9UIiXxEoi7JryEsojZt/My6zOzwAoVtD1a03LNvgK9H6qV/XrKP9nep7tnSS2gooM3yhmCjJXx12+S+TmJMk5fdXS351OeV3ScKzy4LZcsFmNqN7/z7DwyO8XoQUqqHLOp26Dp51nkGJ8CTxsM+h9FBByMnTV2TrjTsOaC/u1tbdFVw7HgaDlpaN53GB5XGZ8W+XK3rHY/rKEJYlQWEg8NwXbV79roXhTQKtfrga3xTc7YT8dDji11nG42TN0Tzl/XGI0qVTFKymE/j81d1DPnnyjJMiY73akJxc8PQf/413RgOCwEf7eyZUS6sW1V43FY3u6iS3pExa6+AojG30Q1EZa4jrNVh2dJ5GSJsKh2KXl9QgZAanN7dBqRoBWqeA3jA6F3Tn8OSMFWRGcLHccLXOSUsXyGkQFQriVuFo8kFEq5w8u8/+mrHTTLzt3avfEtUyVWtfxSPsrGO7oBQOCbC4cU7fj/YdeQDk10uXZu9UFoVwlccEVOfCCpeid6sj5xtronJv1kRds5FSCYJuiP/gkNFP3yNRgvTLl5Qvz1guEspcU2jDIllzkWe8EXk8iEMOAo++J4mlIJQQSIGPbMjeUsEBC0GOJCst66JgmqWcpAXP05Kv8oKnpeHS80gin3LcdXEJj44J7x0ghx20L9HKZVYYAV4UoaIQqzxHpDuacD3PvcX81o5XbtbaWv6A6lmDZyxBXmAvp1x9+DHl1ZxOVnCkDe9GHn9xOKCvLNIU7rvSoyjgy/NLrjYpk06HdydjQmEcprspqSGk23e+lYiEwnoBufX5dLHiV7OEP+SCMy8gkWqbhtVM7aaOtta/kODHAQdHE47uTOgOO0hfYKSpnWHbJYIt7VmLzguy+Zr12Tn64opovuAgzXjkKX4yHPPTYcSjXsCdWNCXGmlzRFFWArhGsWsz/LZQEpUXo80QW5+VbL0D9eNrvAaCnWh4W9tbtUegiivQriMhJJ4ReBQgFV7Ho+8NeK0T8voy4zfzhMdpxsnlFUlWcjVf0793h3DUQ8U++C5QzfHmCoCmGo8BpC+JejFjJLqAi1dnbJbrrRJwu6F5/YIQlFKxVnBWaj5Ocg7XOZOuT9eTTLICqWpcA9lah5vooG2alwhT4NmMtycjnq2XvFxveHx2wdv9h5WyoxFGEynND0cdftgJebzIOc8K1rM1mw8/xf70A/zJCNn3KfbTlxo9dF/puW1o0mUI7Fn7t05jZ82uf74dzHtTXEJdy+V6u6GvfWAgV2mAwkhWacl8nbHKDCWqSeXcKs5/vP/t5/aeXUNcNzfRKAi3fcZWvMatvTEWIeUfAR7587XvSAHYtyD+yEdbCcJ1BHJN1uK2vfYfai3rwF5/xwgoBeSBglGXzjuvYU2JiAKyXkR2cs76ckG5zlgWJZdZyovMcpxuOPA8JqHPwPfoKY9IKZQUrviGcISuraEwsDYF88Iwywou0pLLQnNhDBcSZpFHHkfYyYDwwRHdh3eI746x3QjtKbR0ngotJNaX+N0uKo6bKN9tJcWKeX+bWtQta3wdv9tWBpRDrVMWfA1qmbB59or88VPEckWnKHkgBR90Q97uhcSmiuiXkkJIrmYrXiymYOF+f8C9UQd0Cjqr3K+VW7sRiHtWILAVigrrRbxYa/7tasW/rzJe4LNQIWW7sl8tCFuz2ekKC9ISxB7jwzGH9w6qM3+FlVVNC0FTOc9WtGcBqw35ZkMyXbA+vYDzc4brFW8YzQdxyM/HQ94aDXgQK3qeIbBFVWSmAq1pW2H7zEpUsQvSYaRv8fpr3IGK+Urh8t2r0YlKMW/2IHWRFxyQEO5aowTsMHBnXVI4BSCWPqGvGI06TLoxb3difj9b8e/zDZ9Np7xaZ8zzkjA9IJ4M8AddVNACdhF2O68qCFsEirgfc3j/EEPJlbUky/VuDOCOslULjLrTCt7Xuhz/Qgrm0ueJLhmsEo5Uh3FXEWhLP80h8hCySZir+m0JIdG6Xt9YaxAZ417M3f6Y803Jy/kV8/mYySBESRenoUzBQRjy40GHjzaar0rtXN0vLlh+8ZzRgzsEcYy112HSLM7yb0TiNTI3ILYGiNuCW79T+7Sn3et+ttR1eebmu63SB/v7/boU2CqkXycdXSyYRFtFUsDFKmORluTGWf/NLqr33f6wKqjg9rC3JydiN6lj/7vXWg0iJG4X6TXsu8AK0dRq/F627w4IqLFCd3XUptUrZk3jbtonuYa3fCsDdIRbex52hy5cqWAlsbGPvDNBrJf4CtQgRg67lM9OSc/n5KsN6zTnvCj4Ms/pZDmD1KPnefSVR+hJAilQVboNVrgcawNrY1mUlkWpWRpDphRZGJBFHrofEx2N8O4dEj84JjwaY2OfUjgFxSBcNUMFMgjx+z1kHDVFgGSDGw43HMB8e+0WGckekxA4P5Gfa/JXU64+eQznM4JNzlBr3gwVPx53GEgNZUkN+ZtqwePTV6yKDUf9MQ/HI7qhdBUBTc7W9de+b1sJajEh4YEMKPH57eUVv5ynfFYIZl5IrnyaPN+dn+tzosIH90NFf9znzoMjesMOKlQgrVMA6rtWSmBD4KUhWyWsL65YnZzB+SV30zXv+5K/Hnf463GP98Z9up5CmcIJVVNUgr/qo1lzV84FKV1wq5AOrdA6JaAAMmvJtCXXgtxqcl1SlIaysoSaojDS4vmKQCpCJQgURFISqKCqJGcQDSa6qzMgmoC8ajdb444lKJFSEkuft8KI1w57vBFHPIjW/HKa8MvFhpcvT1huErLkgO69Y/qTHviq4RM1klsdKCyERfqS7jDiyB5ijatrkK4222feVt6uKWzCrUt1WQvBRnpceAGfpxl3vZTjIGIQ+YSbDF8KRFhl2TTRijdkHOx4BzQUGSqKeDAac7HJ+OrqhCcnp8S9t+j5IbZMEUYjKPjRuMd7y5zfLwouc818lXP5hy+I3n1IfDjCsxZlWwLJOFqyxmXz1xH5u3PdGjv2WrCn4yVyhz1U+3SPZdzEgw370fctD59tm3Hthb9lD7XvjURbSWpguim5WOckmgp8S9L2eNT/mh4aZe+Wgbe9APU2vNVW3fKqbVp7O0X95i/+py0G9Bw4RlfgouwY2tCcnmKtrXAkJVi9RQGsXVrOmLqmFHxrrb5Xy2KwwsU5iVDhTfqYaQ+dp3ieZNjvk0+GbJ6dkp9PSWcrkmQNaY4qDIG2BEVBkOZI4cB96qhsa8FYSSkUufTJlSL3PYrAgzBAdkLUsEPnzoTha3cJD0aYbkDuS7RXxTtRKwACowRBP8bvdyD00Mrlxm4zqr4VF8r/YnOCA2tRFgIDYr1h/vQlLz/6BJFkDPKCe1je6US8PepAmVQ4/pJSeFwVJR9eXBAoy6PRkAejPi7SPa+sna03qX3f9i9nSTq0v1KGXK5z/vVizieZ5VxGJMpnC7daMy11vT8srq68RiroDwcc3z9ieDhASoNVplWYaW8ItfBfrlmcnpO8OMG/uOI1XfJfI4+/OhryV0dD3up4zvuRVcGNDUrdnsUvpAOvkQEon1IqMuuQkDMtyLVlWWimWcGsKFnmBYs8Z5FlLPOMzJRYDR4OFTBQgk4Y0A8jhrHPMPCYBB6TMKDj+QTSOqVACQJhkbbySFRFh+oz5qbKosaNX1sCP+StQcRBr8O9Qcrg2Sn/sljz+dmG2XpJkad4PCQY9pGh817UvGALvGwBjVAwGPXACEwJ58UpZVays+ANSdwgjFqKYS4VhpBXRvNJknE3VNztdujnJYO0QEofAtV8ftezdhOnsm49dMG9XpflaMzlxRkfXrzi3qM3iUIfT1VgVbrgYa/LD/oFj5IFZ2XBKpcsvnhC/8lzBq/fI7Sqxklq3cI23qQ9l8e1sRjjYvT3LfX2DGyLtvf19+a+18xn2wT1Ghx6oHP/Xzfsbr5r+29RAVHBMi25WK9ZF4YSD4NH7QNpKxZNkOKNgCfO++YK+1Ti+5rToLqwg0BXd+c8KG4PW4SyzeliY0/UWRPVhf+0CsC23e4+uo0grgUKVgF537Y/pfJD7Cju9VicEiCQoYc/GZCnCasiI1YhYXRMOOlTztak51PWZ+dwOcMmGVlWkBYaoTVCgIeLdm/iDExV7lN54HsQeqhBBzUZER2N6RyNCIcDZCei9CWlkmhlm/g2i0QLQSmBwCOe9PGioMIAqG2AOm3nRh/ft95uzlUGKtAZT0NQWMrpnM2z59jTVwS6ZJIVvBk6GORhqKDcAAYrQ2aF5bP5mi9twc+jEa93YoaeqGqz19bNbbUk6mCdCl9dKowXMC0l/+/zl3ycFLwiIlFhZWm0c9R3JrDtT7rIcCEtvUmfg/sHjI4G4NeA61uarpejxvm3pSFdLLn86gXl6TmDxYK30fzNIOT/un/IG/2QkW+h2LjYBl3n7+9h1FeC30qFVT65jF1AaVrwPE15stjwMsl5uSm4zC2LEjbCdZdZSwbk+JQopGHrASgtItd4qw2RTAiFpQsceh4P4ojjwONBN+KNQcz9OKDrhQS+RukCVUPe2loQt2jBlFBYsCU9L+CDUcCD6D6vPTvhH6YLPtosOH1Rcp4ZRm88ID4c4sW+gxNur3+9V6tH2hl0OLx7hNaai5MzTF7znTpds/U8beuB1Oe3QoD0KK1ioywvSsvvN4YHKdwJ+0TZEi81CCEhkLtMacezVNEGuGejAGsIPMFx1OVB74Bfzp/zdLmhF3QZKQm2qlYZSl4fDnhvWfDF1ZRpBsvpjMXTZySnj5hMDqvoqj2F1gJVEPPWY9J+z0kzaw0NiNUeopBLojAYTAPS1H5yTUnpZqYtAVynzlmzzduXVLDSX2NgUwtfs3UaodBWsMkK5uuMRRP1ryrhf3NPwoqdEkLGRTiyDURwA6kVFSFwXlJBBXfcyvJodOstzkEToF4bqg0SaLVWwmWVKSVt8L8VgN0mrHCVxv7Uz+PcUvI7EP7A7kZq/qxxsEF7An/Uw09HpGlGukwRQKA8gijC63cIj0aYxZpylZKtVhSrBLtJsMY4L2grzsGlTSm8OCbodhwwyqCLN+igehGyE2NCn1K5AD+3mSrLv2I2RgkIPLxhl3g8QASBi5JubRCnQNmdDbsrlysX17eIteDusqsAOtvL4uUF09Mzli9PUZuMbmE4NCXvdjo86EYoNGiNFQorPc4WG35/ckohJa9NxkziAEVV5rft6GgnOe9MumYECqTHRsPTZcK/XM55riMWKiBTnit+U7kIdx0JLaEhqqMGYfC7AZPjCaPDIV6oKjN1W6ClZgd1ppouSzazBbPnL9EnrzhYr3jfg/9jOODvjse8GSt6osQrcicwzZaBNSuoKqEvPUrhkxvJJjU8Xq94utrw1SbhWZHzsjBMjeTSSFZWkUpFLjznUZFQSnfc5cLI3Thlo7BqpAUlLMpoAm3o5YYjrRlScLhIuHepjvlJpgAAIABJREFUeD30ediNea0TcLcbMAg6+LJAGVVVGqyjsnFrZgyUGkVJrDR3Ip//87UDok7IcLrkV6uUF+fnLCRoo+kejQg6UQW5sHUVmtZjVr6kO+hwZI7INimr+dLphUAT7LhD5qL1XiUkrABpSTHMTMjTVPPRdM17d0ZEwscrCgJlHDZABRHbCI6bEtFrq8KWSJMzihVvHk34p9UrPj454dC/y2AUIEW1Trrgfhzyfjfkw6nhpNSsS8vm5Iz0xStUp49XH7U0fddn4rLlCdifrN3+3LDXm/S5Vkr01vjad7Jf58lbzlbb2G0+88d4S6UQV+BEBkVaWGarnNkqI9cWIyWG7cNuh5hvUQi2GQE7rXkOe9d2Profs3dd6uwWY2p/vvYQisprIOz/9gA0rRY9t69HG1d6Bz54T9P/ptqOKGqQMyqcgkqTbpitcLy3lAIVRwTjIeEmI80vya2pAoMFMvQJ+l3sYUmY5wSbDL3ZYLMNpjQVUFWdDy+QUiGVwgtD/DhGRSEiChCRh1WuAIiW0uWNs+sFsaIK/vM91KBH52iC6HQwvoepAwCFaLZtrb2KGxnCn6cpnJEsVwnp8xOSF6/wsoJhqXkoBO92Iu7HEZgK9U965EZwsU54vpwzCLvcn4zoBRLKrDoiaFl37WZ3uIW7JBVGKl5tCn51MeejzHAuAxIZUAqPxshqJLjY7a+uCS4MXqA4PJ4wORgTdyKk2mWWdQyLM8IkJi/ZzFYsXp5SvnjJvfWKHweSvxv3+NujAW/2QgK9QZZ5ZUXvpjJZIZ3wVwFaeCy14DS1PF+nvFxt+CTJeZJmnJQFU2FYSEWuPNLARyv3Y6SHta4uh1HOWnMDrN2rbp7G6MqAsqA1stRMS82lFoRlQacsGKQ5E5HzYJ7xKPZ4qx/z5iDmta7PHa+LLzXSFIiyAMqtFmRcWqcw4CvNw26A8gaMIp/+6ZRfLJY8P9OsrUPN7N89xg9VBUro1mPr66mzLxR92eM4O6bQJclyA2XLAmwTwQ5RtN1/hkJKVsrntDR8tkr5op/T8XxiNF5uUco6L4CAbcxJ+x57HgKjQW8IVcRk3OP4bMzT9ZxXqy4P+wfEnueOsHTByAt5q+fzfhTyWWa5LCE9nVJ8dYI9uIOnbfN8tgHTTgAJ0YjfazTfvtDg+dsdn4p7ry3Eq4/U9su2NG9lOKCcv8jWaXL1fE3DuPbTCbcw5S2aroL2LIrcKKZJxlVSsMwNRRX1X1vgtQ5c+zmuGTzXtPbtfbcgQ6L2O1QGUr1mbe9avSJbA8pW6369VesPVmwVgO+lEvCdKQA3WaI3topybKWAN0hX2282Pf5Hm23/1FqgqUGKRKMsbtEHnSJgAOEpvF6H3uEENjmlNhSmdG4p4awCESk8QgLbw9VXN+gqP1pUQZGm8grKGmRDOteVrt5z+a9iu16N4iuazWiURHZiosmI6GDi4gekdFjU+3Nuoii/uXX8n201xgJsPXK+MeirGcXT55izC1ReMtAlb8UBb3Yjhr4EbZ31rwLmSc75Zk2h4M3xEcNuRCAr0Jv94Kb91qap6ux/YyRPlmv+6XLJcxmzrND+bDs1rlEC9pUnd90LFL1xjzv3jun1Y6SyW0O9WWfRlPW1hSGZrli8eEXx8oTD1YK/jH3++2Gfvzno8ShWUK6dUtMGM6oikK0SoHy09MmM4iQp+HKV8/tFxofLnCep5hWSmadIo5DCV5jAR/g+eD5SeSglXTaAdZHUWkKJwWgHIGBsdRxmLcJ6jey02qK1xmhLUUqE1khd4JsSvyz4NCs4SFNeW6W8t0j4YNDhJ72IO7HPOAiJgkrIlQXCVnOztkrd1EDJ/aBDb9KjLwWaGf+43PD01SuW2sWAjI8miMgDtUfFomLkCvxIcXT3kCTZoAtNts7Ywfy41RNZK/0WoyFTipn1ONGa301XjA/7jKRPVOZEaYHwAmeK1srTNX7fNmQ0lBnCF4RhzDtH93iRfcZ5smaxGRCNOqBd2mDoZTyIFT8Z9/gfJ1PCXJNdrShenJPdvyIoLNK25rN/u0YP/hqjq/IY7PexVat20ym3onH/8/WB0d5KVsy8EdAVrkD7WHDnb/5/9t77S7Lkuu/8hHkuXZmuajcOmMEMBgQIUKRAaWV+kXR29w/YP1faPdo94opLUaIgOGIAjOtpWyZ9PhNmf4h4JrOqzUAkMDxS9MmuNM9ExLtxXdz7vcHyN16zrBwX25rrylGicUIH67/z6vle4Wh7PeBvPjLxG6MfPKJWUZAMyWFwwMBD0CMctuNvsQBuoaN4+v/EAeha4KCv3Mc/NHFjOk1IGWvzuV8y4b9DbzrLfv/b7m9QNFvNONRg94ATAp2m5EdHyMazMAbrt7im6YA4AIwP0f5CCRQqXrUNIukXU7+jGQjPDgEobt3GbhUFic8yipMjRmeniHFBM2SIB9O0p8/uKQK/x9bm0sYcauE8qvEsHj2hfPwEsVyRNoaZrfjo6IjzQqNFDCaTGisSniyvebpYMMlSvv/wPoUmCI8Ooe4lHoC+E+GlUrzOeb4y/GpR8qvSc5GM2ckkVmY4aMMJHNCoSATFdMT9t+4yno5QieytLx+Y7KBKO94I6vWO5aMnmK8ec3ez5Iep4H97cMqP70x4kHiod/sKjRAxriOm8iUJO6GYN4KvFiX/75ML/utyy28NfCVTFsmYXZrS5AlilASvVZ6RpClCKaTwqA6FO6TZGW9prMXEF9b2ACtO9LItAUjBg7USbx3eNJTGgDGsa8PSNFzaii/nO35xveS/pZo/O53x/fMj3jrKmWoV6lXYGvwQqVCEbAG3YZbk/OhsBnoEn38Fq5LPn7/gyjSheuGdY0TeIte0z6Zl/kGhToqEswdnVGVJXdf4Js6nUzcJ5LbtLyFpgJ1UXFjJzxdr3poV3Cs0RxiyskZkArJBH/YuO/zQ/hi8Hnnq+fj+XX71/HMWqxVPV0ecHh+TyLorFXyap3x0Oubk8VPGZcVWSbbPr1l8/oQszdvQk249+0Ea5p69LYb3H/auDYS7uVj2MjoHFpOAQZbBwTkE7uQHYw9Lfl8VPpyf/jaCxitKq7hc75hvDTsrsKho1Awscj9Ykoc2TVt8pEu2vckThud1U+DtLcdFpb0T/tB5Afbk0XDCgm4i5GtwcP6A7feIAzDgnC3MI4ckJ2irK7VT2hvfPUDK77xF7ff+xPvdpjn7W4kkjCIAE8kYbeuyhPTOEVPbsBEXmOUG6hrlXAB6EwPDMV7P7V1cHMyO4Da30nDfTSBwIgQkkiXkd44ozk9Q0xFGqu4SA1ZDC6T8+7f391tf/rPPVZbO47cll599ye7FnLw23PGWt5Xkg0nGceIi7K8FmbMxjserJbvdmu8cHfHdWUFq111U+UEe0y2diP9JiU9SSlJ+dr3iJ/OaKzFiLbNQHCYqaS9VIkLnQXjyIuP0/JjT8xNUouJ+dKTXSAQtM3XG0mx3XH/5BP/0BQ+3a/5RLvlfH5zxL86PmakGmgpMm9Ovuht6oYLVr0Lp409WFX95seJvrlZ8Ujme+YJ5FspDN/kYOc4pRjm6SNCpRiqFkz3KZcd6hUN4j/agEw0kVNZincWaoAxY47HGRWttULlPOqT0kIStBIzCVJq10dSNZt1oLuuaR03NL18s+cG25J+cTfmz8yPO0jRkDVgfLf920QSPD6IhFZIfzcb4B2ek8pr/sNrx68s5z+VnnPE+o7NjVKY750wf3BY9Z8IxmY05uXdKVdWsLpYEkKMDvtQVZIgf97L6BA2SBZIvUPxyU/Ge1jzQCRNbIcsa0pSOcwkflDRPUFwP7xO3FhMsD0cJ384KPtte8tV2xbtVw4nWQAPWUCSa+6OUD9KCR8ayqmp2T695kT3i/tvv4o3vjRTRv/qhePa3JvZbW1cgQKz31obwgbw9vXOjc3Lwcng3EY02ge3o7Nbj+h7gopHnkBgkpYerreHFqmZtBCYCAQ2v9fIQQDqPaS/428CpyMW9CBkULsQfWW672KGEarcmhrrGDYzEvbP/nnDr/87aH6AYUK/tdeT4EokellJLwvvEu2fJvsG92/t3ez/Dp+h7xWPv5u3boQY83KsSAi8FLs/Iz0+RQrFNr6jmC9yujNlZYUuh6/1ACfEH8yEQ/QJ7yZx0wX9aQpEzvnNEfvcMPZvgEhUXvuCQJtt82ED+v3+ivG08gpAgqpqG5npO9eQ5LLaMGs9dBB8eTbk3Tsml7SL7nZI8W1U8rWryNOd7R6eMtUDW0UMwuHpog7H6wW8CkBqnUr7cNPx8teO3tWWlRlQiCRkVYnCpG1Pmu991ljA9mXF855g0TeLW+W33DfK82VYsv3pK8+Qxd3ZLflhI/tXZjH92/5iZciHYz9S9JQIgJF5FlEKZcLGz/ORqyX9arPnrVc1nTnGpR2yTFDPKYZKTjgqSLEemAqFE2IoWPmBDRAnhfKzSJlxUUmIpYEALFbxWSUgZs8ZiGh89BCZWAvQgBF61hboiSp5MsNaxaxqqRrHWmus6Y25rrrY1z59d8XS3489Px3zrKGeqc7SVIchxuDaNQSLIleCPTsZUUiHUguZiyWeX1yyKZ6AU49MjZNoy56heDuS7SiSzkym73Y7tdoPdxMBNfwumw/BZu+gC92CEZCcTLjR8sqn5bpbx7WnKTKeoukY0DiEFqAGC4lCoDi1UDziPsBbtGz68c4en5YYnZcWj9ZqjszHKAs4gnWGSFPz4rXv89tEFl8byYrVh9eQFqVOYnYkRkD2P7NCJD2n2gHP2jjLf8Y42bmjP1r6ZK/fS1hlvkZ7aLS8GcQY3rhFhwg2SCsmycjxfVSwaR+MlPeRRr9kMjZxDaSD23g2EdMcHb0Ibd9+Jw2sJpL8ZUB3e3OKe7VhD7Nn/6DEAfiBD9301t7TWNbz3XWRcQFsdcJiG8oZ92NOMbxJMhOW9pWt98FwvEVoN00HA7x+NSO+EgCwhJdV8jisrsB7heqa6p7X6YX/6MD1/m/s6LhArBV4nqPGI9OSI0fkxejbBZ0lQRmS/wPuAoDdp4nf3rPwOTXhi7r8lKWu2T59hn1+j1zvGjeFcOL57MmOaKRQ1eBMsdjxfrdZcVzXnRcH7J8coW9NVt3vtIFpLSYJIsF7zyXzFJ7uGZ16xVQpz255La14OP4uQIjWejjg+mTGejkCJCFe7ryhCINymbFhfLlk9fsJkccWHGv7pyYR/fDblPAGamAe+ZzkIvNI4nbERCV+ua/7L8yX/abnh56XhU6+4TgpMUSDGBcm4QBYpIk/QUsXF0q6fyItiSk1robnoWWsD68EH97yIaJxKoZREJh5pJNJIrDFY63HG7S8nJfFC45UHLXBJqLRXK4etNVUjWJcVc7Plqqz5sT3h41nG/SyLWwIe0aIZemIxI88sUfzRNMd7z7aq2awqnr24YJWlqFSTH08RA8bQFngJ8K2evEg5Op6wXk5YVAt8Y7v57R8WB6yhF4MeQSMVayl40uz4vGp4Oko5S0akxpBUDqUC8FLn7hkaD9212+9dUHjMlgd3ZhzNR3y13PDoes737oyRorVWHbny/PDsmL98dsEXpWFRNWwWS64MmLKJnq89q2ZvaL4riNS6CFpzYPAdByghUYqL9tg3FGHDa7T3EG365V7rzZHWR9EgWTee603DctdQu2FC+H4qYhsDddivflytWSUGYmegjHT+gf0IiBsyICoyw/HtG4PtiG/ynr3whG9g+3tXAHwoIP7aowKX8VFbummjBubVu4+HqJtv1ES/BgM8rhxY5K/pn2CgmOwXwUQEl75RAj0ekWmFTBU61dTLJc1mi61rnAmxAN6DGgj4oVEAdDDr0CscneKjBD7N0JMx2ekx+dkxyXSE0ylWqqj/t70Lwv/NpujrTuaw3XbeLQth6PogQuk4T2ocer1h/umXmMslxa5m2jTcywUfnUwYJRasCecLiasszxYLdlXD0eyU88kY6rK3/oe3fhn2AALQOJmwqT2/vFrzWQ1XIuyph9DyIbhO/G+IDIUH4dCZ5ujkiKOTGWmmAxP2oieXtn6FEFjj2M3XrJ+8QF1c866v+KenR/yTsynvjROot8Htb11/T2So56AzVqR8ujb8hyfX/N8XG36N5EUyYplm2FFONsnJpgUyS/BKhiDB1iLsLzf4Lq4mD164yAb7tScjgXoRIl+kBK0EQulQl94qrHHUlcE511Viw8d9aAUoCSoBrfHKsUsSmlqzrRPmzY6n1xUv3IJlPebHp2MejgqkcPimQfhBTIdrgC3nScGPZhn+wQlP6gs2qyWrp4pVnqKKjETpG+TXriKtBdPZiPPzE8rFlsrUPVJcK5xaRa+TGO2kBcXCyBALcGlqPqsaPqsMD4sxuSqZ1TU+8Yik7YO5nfxaxuM9eAumZDqecTIe8eh6ybPlnKY6R2mJ8BK8IxWOb09S3k/gFzvHE2dYlSXbysW84NbMGr7aCWjHI/uxiUOrTHRIgrLNNqIF8TkUka9vfjBvshOOsqO3XjhH1k9Aq6yMYLGtud5UlAaGYMei85YO+CIDE2eg/PdgQC9TXPa/bNGl94W/6B9Tu2W2hyDar6MwpJvzI/5HVwBuNH/bhzex2uT+5zeY1oNlMDh3gIV9oLmFPf597fn2a7dE6Lun7JVA5wm5PmY0ytktRmyv5pTLDaasQoCgtWgvQwxBS9CiB7R0PnrzWoVFhAI/QitElpIdzSjuHJMdH+FHecQGkB0Qa68tx/rUr5qnSMj//Yb/vrX62qN8UKOkA91Y/PWS+W8+x652pLXjyDve1pL3JgmZa4JwFwExsVyWrDZrchRH6ShYsmUVheYbrjURhFLtUx4vdvxmWfLcatYqx4jk5hD6KWUvxUsEwJnZnSn5JMdHC0yKFl88prI6wHmq5ZrdsxfI5xe8bQ3/dJLzL8+P+fYkDwBHTbVv+QsBKoUkZ+NTPlnV/PvHV/yfz+Z8KjNe5AXVaISYTMiPx2SFQiY9TkTPfPeV5j5L2iMVCCnQSUKWpHjjaSqDMfbGWu1WqxJopRA6bA9opTGNoWksjWmx4AfWtZKgRIy5sDSpxpSKspRUIqNabliUNdvK8K/fOuduUSCdiLDBg20dE+KpT5KCf3x3xhfbmvWTC342v6Z8mrMZFRzpEA/Qby/uP8osSzk5PWZ1Z8lldUlTWgIbvCFO+mfgBV2ev5QY6dhKzeOy5jfbmm/PphzpjHHTIGuP0A5yxZ4C0ArgQ55nHfjg4TrOxxRFzrLaslysSe5M0TIAPinbME4s7+YZ5xtLbi1SemyHPzAYAoPv4vfitsl46VKNUfq9Y+BVB996wT4l0Xfhr/scuZe24ViF9Yr1zjJfVSx3NY3PBkfvC//wpWiXYbzpgVDvFLhb2iGruPWwKHdaQ83v90a0ikHMlLnNaHXwP5EAXymtOwIWrzxS+mhc+YBr/0aObdHmdt7Sn94nNPjbxgF8DYt4KKwBKxUkAiULklQznU7J11vK1Zrdco2rKmgc3li8MyG3GmIaVqsRO5wMlh9JgipSsvGYbDYjmU2QowyXJBEbQAzwrnvPQtc93y+ev18f/+uVuZ7F+pj6B3JTUT25wn/6GNYVmfXcFZJv5SkniUfVMaBLZFRe82h+RWNL3j4+5Z3ZNAgFCz0q3uvGKfBS41XCshH85+cLPreCucioZIq9xYLsT23T1QAJKlUcnx+TTzOEiiL1oJZEZKWYsmb9/AX22VPulmv+JNf8m7fO+PYkIbVV2PN3gxx/AV4rUClbkfGz+ZZ/9/SK/+tyzW9UziorMOMJ+dGU7GiCyMFri5U2Rkq3+9AtLfc4EFIIpIQ8z5hOR0ymBcfHJ5wcnbC4XPDoyycslltwoZqZ9RaBCPUBaGGsA70JCVmqSbQk1Y66tpR1gzP2ZmS5AoQOKH7SY4TgmhonoDYNq4uKhb3g/3j3PqdJSqJtyNv3pmP2LZpPkcL//t49Fus1u/mGX11dcKUUo3GOlGOElih5C1cRkKYJdx+cs17tMLZiv17rUEBB58rfaxKrFJfW8VnT8GVV806aUDcKXdegHGQZEAGCboWkHdzPW6grzscj7own/Ha74jcXC0YnM6ZaBa+QCwWfvn085f7GMN44UuvYteELt8qYgSfVi5sBacPnszdFLT9u+Ykf1reE29IO2zm7pVkcIcyuVQoHiA1xOVkku9pxvdqw3DYYJzt8wtCT1lMl+iUygGsdjuwQqqjzBoh+PH1/h8GgB22gAYnBaaEfHi9sKAiJ6Oqx7JUHfmmu+zen/b0rAALr+9u8RgC9lHH7Lvitv+4btE7h7JGZgjI7iModxGcEgpI98fge0/pgUIPOBIJsgTFCP2XIMFKA1ugsZzKbUpzWuLLCVTWurDF1RdPUeGujrhniB4QEoRNUnqGLHD3KSYoC0gwXoYBdRAUMozjwZAjCnpW/2e0wzUNF4RVa8msn97/jHO+R3uE3O3ZPLvHzFapqGDnHgyLhg5MjdCwr65F4qdmV8OnlJcpa3pmMuT8ZBXAga+nq2u/tyx32M/4mFbVXXJSGnyw2PHcZK5VQoTqPzk0LYbD6hUcmmuJ4zCy6/ofrPsbFRfrz0DjWF3Pq5xdM10s+SuCf3zvhg+MxE1kjbZvn394r7Pl7lbAl4acXa/79szl/sdzxidRcpjl6OqU4PiEZ54hU4pQLTKg3h2jp2/sAT6wVpKliOprw4ME59x/c4+zslOPjKePxGK1SPvvNI3bbGoTGO4+xBmPCqzaGxhmsi8pEt3Q8SghkkqBkwBaoqpom4gT0fXHBGyAlyASEoJGaRSkxTUNtatzVjsI+5V+9fc5bo5wkISoB0HlfnEHZitMs4395cMJz57hcbvjqxXNWj6dI/RbJtDh4+nFbB5CJYnIUgjab3TVVM5j7w9Yuq6HxCjRCsJSKx43h0/WWPz6dUaJIHcjGIWoPhQoW/g06bElxIHyd4ayY8XAy5vEzz6fX13xQP2ScyBBSEGsIvD0b89bVhqNtSeYcVavw3Sa/bnzhA3G2kKoxh66DxfB0VUNb/aezcLGD9EJ/29UHLfDbNre/+/9QzvrwRBsnqZ3kcrVmsTWURuBIcC0qI20fBuMYeC9frl6J/Xftf3ssQdw49kbr7KeoDEToYC98jC9h8Dz93mnC40XzzVUEfo9bAK02ddgisYi9I4E4nQMr/mugBx9cvQ9F6fRF7+L1g+tYdgT68me1LzgHrVMogzXuhOjqxgshUcqjsgw98mAs1AYagzENxhh83L8WiBD4IwVSKUSaINMEmWiE1lihsMKHoj+tEt5a/y2PHbjFXu1TuW0Ab958ZMivcyrs1QAQ4Zz2rXSOerVh+ewF7BrSpmGM5UGe8d5s0uf1y1D4Z21qHpUrChWK0BRaQN3QWxYc6DMD60tAR2tSs3Dw603FryvDQo6phOwR8Nr84RvT4rqJTTPN6dkJo3GB1rGeQHwOQTjG2beWertj+fwCNV/y0Fr+7GTMn98/4TixaNMMahf4rn9e56x9wm/mFf/+6Zz/uCz5xAvmRY4/mpDPpqTjDJkonHR44Tr41F4pDZqIkI5ilHJyZ8bDB/e4d/+c+/fPOTs5YToZk2UpSqc467h8fklRpORZAoB1SfACWEtd11RNeBlj8XbIegMz9FogpEYpKGtDVTe9EtB6IyRdEKaQCY2QrGQdrL3aoq42pFnOP78/491xEXwZpu5oB+8QxpCILR8dT/izsuarqmK9W7J68pTk6IhxnqBVcvAIwzMRUpGkiqPjY9bXJdVmfWAVMhAy7XetVhdoxEjYSsmFs3y53XF9MuVcaQqv0dagqgbyET22wW1CMz4rD1hPkQruZCnHScLjcsdFUzPzOYUQ4A3YhqM85+4o53TZkNUW5du04j4+6rUt0vdQVLWCvt3tD9BAcVtS0BXPuR3kqB3NgbItBlPY3Wlwuiek/XnJsoLrjWHdiID21wXixlF1SliL8im7a9+c1WGM/9AiH3wcsAURhXcPVHTr8OLTGnpqhzQy4BuDtpeY9A1sv8cgwAO3EtALrm46h7/E84Om1RL5MHrzda2zi7tn01NAj+3vEMIhRbt84r75a24huv77aDDG64r22iHgRorgA3F4hBaINEFlIJxHe4dyB27rFhcgCnkrQmnSLhob2cUI7E3hzZmNl3zFQG4opvvH7hfwEf3/B5e8aSz7GwcMkblDPrFDNJZysWH57BIaR+4cxxLuFilnRRoq/1lAKSovuKgNF97wcTJikuhQP93ZWxde37N2BUahKCReKq5Kyy9XG56gWCuFU2362uBae96EnvEJLcnGOScnRyQ6CVH/YsAUOiECpjKsL+dUF3Pu7io+zBL+5HjCu+MkVvRr4hjCVliA9k3ZkvLl1vAXTxf8xfWOX3nFZZ7ipmOK4xnZOEckIiiwg7kVTsadrNDfNEs4mk259/CMt997iw++9Q53zmaMxiMyrdGDMTYurAUhQiCYEAKpgjjwHpIkIW1S0rqmrmuausZah7ft2g1KgFICqZIYtOvDcW24th+sYyUQIgIQCdh4yxPnoIHicsUkVYzUhLt5Dt7EHZhIW85Cs+MoT/mj4wlfbUuePbnkp9dXbK6uSGYFOgs1DgaUGddXeMaT2YTxdMx6sQupdEIOFMbblP2WNoJAqpRibizP6oZnTcNbWjH1CWmrAFhPh6Q3lHxDodGmITqHcA1TLTkvRvyi3PFkW3JvkpIrGdaUMyQp3CkyztIdRWXQzmF8VHQ6a/2QgfneUNiTh6Ibp4/PJtgfIXak04Nbntvytpfa3L5b6+0w3Y112W5Fhbgl4yXbBq43FYvKU3mFFSGdWe6hwNLNfeiK7wyuVjl4tYEYac8Pn+swNoGOiR6mCPY/tRklLbfd5wtvHIP0DWp/gCBAcZNuhj/T6QMQ3/cxFH7w/xvcqnv5fu0eHNCxzrg2eoMxoIjd1kTbsZfdbyDMfSQY1219ux3uAAAgAElEQVQgxbLCMliJzqsorAOmAFEDdwLskKBu7F/F794gYPHV7Ta160D4337IG122fZRdvK+XKO9ILMiyob5esLu4QjeWsXXcSzR388D0qCx4gfeKVWN5vNmyFYKz2ZRJrgFDF77b9e2GGrQ/AKWxXnK5LfnVYselSNkpFUCVOo1xIPi7eYgWuvCkRcbkZMJkOkKpnhEE2hUdIThjKFcbFl89IVuteFt4fng84Xunk6DcNFXMe49KipSgM4zMebq1/OWzBf/2xYK/FTnP0ox6MiI/nlLMxqCJqbE3lS3wSCXIMs1bD875+OMP+OCD97hz7w6TSYEUBikIUEceEBLvY2lh4SNOTWR57boQkiRJSJKELMtomoayLKmrmqqqAyaAD3Sj8DghyFKFkAlSeerShurFbXfjXFvnIQlli43wLJ1DoPmbcs3Jsytyb/jn750xTlKEr4ML27tgCRoJzZZvjSf8+dkxX8yXPNqULJ5dUM2mjEYFMlM3t2KFAAVZkTM7mbFebliUVyB07KDsGdGwv3vCSAUvgLBcWMejzYb3TydMUeSx/DdVDdnLqki2zREepgfbMNWKe0czzPyKrxZr3j8ec2ekwTcxPdRynqc8zDWz5Za5LaiVCLxChPm3roUak5EkLB0uwvDVDSnk6u9z12E+UXjn/L4nI5hlcjA3Acqnn6YBfwLaDf+Wt1gUuwau1zXPl1u2Fqwf4vwfKDLt+j5Y5wdqwl7z3nfBercJgXaMXUD2K64VDu2VIWi3A77hZv4r2h+gGqDgZbnpHV12WuSQSn+HSRZ9gQcnbG+FDjSMEFIYS5+6Vy/V17VD3ebW+AE8A12gs+Bb760gBo3L8GOHmf+acXbXe10fb2xxtCQv3yhGMHqVbxhIvs2UelUnfADEVc6TWY9fbTDPLxAX1+i6ZGx2nBU5x7kGYWNkv8Kj2FQlz5cLtJDcOxozTYjogO0Nhy5DCIu0jZBq4wMCit66tjzbVjwuDRs1plIyellu7TRDSDghHKNRyvHxBKXBS3tDwLQbTk1l2c2X1JcvuFfv+MHxER+fTjjKBFTbCPbThjkpUBk+yZlXnp9cbPh3zzf8QhRc5Bl+OqE4nZBP81DJdjj3wkcA3fAAdKo4Opny/vtv84MffMzbb91lPCtQWiNkANqJmyGdteOFv2VV7gPktONKlEQKhVKKPMupyjooA3WNtRH9Le6TJkoi05REWsqdwRgXvXktWI/vF36u8T5nScVTn/LX5ZbkYs54nPDj8xGZThBtsKSLz7SpSHXKO6OMf3HvnF9+dsnPFgt2Ly4ophPG5xntHW8AvEiYTEdMjkYsrq5CsJ1QdNsoHSkNhEf3qENefSMcSxo+Wc757smIEwkz4fHWIXYlJGOQLZs1vJKPOcsoUdydTCik5mK1YbNr8JmmyyBwhrtZynu55g6WSzwbH5HsZET06y7YRqfLMNiO7/UagPAC70QsMBn4jfMiZBXFKVAeAqJle2q7Jmyki4AyaDE4kptK6dBn4IOSYFFUHua7msv1hnVjMSSRE7mOLYl4drDy45oemPoi9s9zEOPoW13YYp3H2oEXphu+6K7SqtJd1sO+zUkvt/bvfTDMf3DtD6YACL+vGQ925/c+D8+67f3L2r764GPUpgspcy1xdJQQi6HcYmS//J7+5rcHlvJNYXtw7kGef+A5vXYw1EZvuNVv6ai4+dVrmj/43x/82vZz+JM/GLrv1tX+2AbXbnPh8aGcrIfEeerlmupyjtiUpI1l6hseFlPuFElnGXs0OM96W3K13DCSOUURLW9bBUuwy67ye/260aTEqYwnmy1frHZce8lOaWwHzXo4jmELDE+lCaPpiPG0AOn2T2vv7QI2frXasL28Zlw2vK/gH52MeG+aoiPEa4f0J9qMj4ySlJ9fLfiPV2v+1khe5AXNbER2PCGZ5gglo8IRrKsODEUE932epzx86y7f+ejbfPjdD7h3fkxRpEgdrRy/v+rauIVbZ2wvQGooAAVSShKZoJRCa02SJJRlya7cUdd1N4dCgNYSKQVSSMqyoW5MD+DSerEEoBUUKc7Bwhs+rzTZrubkyQveze9xv9BkytMXewqeANGUnOqCH56d8v3LDRebmhdX12xPTiiOjgKXa/EPRE8qXkBaJIxnBUmR0Kzqfrg3jA/fP2TXa7tOKbZO8lVleFZbHiRwJhVOSlQdEfpkK7jU4JrD2bahg86ilCLNC06yKau6ptzV+EmBlzoUTXKG0zTn3UzzQEq+tA6tPE2LPigU7ZZNv04PnmwrXOM8HvKWVj0Lcj9uYQx63YN403mKupkSNwO29wWtDLgpSJa14XpXsawsBh2hfkW8Q3+Fbrb2aHegz/ibLnsYqP5+r4ft4PfH7Ok9zW3A4YFAEHueQbrdna6H3n9dBvwHb28KE/d31KIW5WVLRS89qm1hTtvQlO7bN7pbeNy+I8ohPnt4hoP38XcnPV7un/Pyu90k868Hl3Fw8sGVb9zX0ycw+P3vutdN2n7NTaMChIjWQ8DldsJFpallBSEiv9tnjK/QBx9gTZ2PzKSFJBqo8a3K5YOlqa2nWqzYXS+QdU1uDEfecj9TnGaqD4wTAmc826pi4WqOJickWRESQfdy5oeafdvfg+mTCidTHu9qPtuVLIWgkjIU/Wm1MB+T6GPufs9JwwSPJgXTowlZnnRG1Q0fjwdT1uzmK8z1kjPn+NHRhO8eFZx0nos+oDC4pBMalfPrVcn/d73mJzvDM52yK0booyl6FtzZTrVxIcGxawmKrZCeYpTy7fff5od/8kf88Q+/y1tvnzGeZGg9QHkUYWsr7M/LyJDFoMTqYErFwW5ox+d6ApQybA1kecZoPGI8HpHlaR/5IzxSeBIpyRJFnmmSpHVhHFC5FGE7YJRQFxlXacanKP56WfKXTy6Y26DAIZKBRQuYhswbzgrNj++e8i0N2WZNOZ+zXa/j9kRLxQMrWYBKFKNxwex4EsMFhoJ/uOAYMPiWjwmcEFQiFAn6qjQsnMCoFCcU3oBv2nRIFYklWrBDAd3SbIwHSpKEu9MjDI7trqQ2DnQIysQZCuk4TzUPtGLkLdrHkDgRLf19jT0IU+/2vvPOY40NUM7hizAzvheTzoP1LYy56PPdoyIkUHQxDD6U7/Ve4r0Ic07LI8K6cj5485zXVEYwXzUsto7Kqvhb2/d2jsTe9YmwwkOI4fBqAZNEz5d8mzouu3iGdpy3KURd+E87AbeY977jgW2CYlSHvEP62wWaEMIL8c0tBvR7VgBg6H7ab71+OZyt9mFLL6Mn7uvNZV8co635PNAt/YG22wqrLrf2NUMYDCX6NQ7+0TONPaSIl1zY778EgSDF3rnsA34ddOV1Xb/Z9/5DG8DYEblvC8R4EhvyjlPrSIxDW0diPYkJ32XGk1qPdhHfv+v3oOO+Tx+TxlFdz9ldzZHGkVvLsfDcTTVHWgYPAB6koDKGTVPSaDg7PiHRaT9fh2Mbakbd3zgzSlN6eFrVPKkMGyQN0b1ISyi3PZDws5CSydGYyWSEkjehk1t55r2jXG+prhekmx0PpeBHp0c8KBIyb8LYBgqLVwp0SuUV//liwd+sSz73glWaISYF2Wwc9rK1x6peMXUiMiXhyTLFO+8+5I9/9Ed8/L0PuHv/DkkqXlIXKQb2ddTSU81w+C2jf20ToBNFlqdRCRiTZ2lw/w+urqUgTTVpqgOi4G1WgIhKQJ5R5jkXScZvLPw/F3M+31p2PgngSEIHa1d4wIKryYThT86P+XiUcmIamvmCxeUVzsYCRn642sO9hIK8SDg6miISNaCh9hh/KE8ZPniPoBaSJZpnZc3KShqVYtDhKi20cztRh2ZCd91YDdE7tJI8mJ2QaNhUJdvGgIxKk7MoZ5hpwf0ipcCS3LJ9E57dkO+4vbXonKOqapx1OOdx3mOtx3qBdQJrJcYJjPUYI7BO4nyIn7FOht+twlmFsxLrNN6nOJeEz1bgTLiOcwJrFcZpGqepnWa5MSzWDZvKY5zGe9VbWw76wj0C4STCBWEvbXiJECTVHzt8DSoiSR/O7eb5hrY+IGIO1//+Y9rfYAkeQU8IbBF+6BcZPoRvdnzAH2AL4FVtINFaw5EYkdpaStx8Rq9q7T58G6nv9stkDbTUAdJZvI+IPqbfKbjzpeeIW63GVhnpjxpcxB9+H7/+HfXKmyAZfu+ewocIXAkoa0gcJIZQnMSHynDOuY7AhaTDQPc65OwbJWmkoBnyORH4qXICWRrM82vM1ZLcCXLnuZuk3NUJE0G3x+ulYlVvWJc7cqV5eHxEqgQdROwN7rw/0m7WpMYrzVVjeFw1XBhHpQR2L0j84HoH7hSZakaTEVmRdle/YSx4gTOO7fUcO59zzzR8WKR8d1pwJB3YElxNCGm3YX9YZ9Qi49mq5K8vVvy6EVykKc04JT8ZoQuFUxZ3mO0Q6ShLEx7cP+Mf//mf8OFH32I6K+hwEYbT0LVgjXrckOqHYu+WOdy/p79l3qWUpGmKUiE+YLvdUlUVzrnO8EqkwCcKnKa0NcYOJrC9pJSILMHZlJ1peGpS/mu544+uNpylKe/naSBGZ8AbWgUgcTXvTyb8YDbm57uar1YL5s+ecnb/DKnSIPDbehHdPT1JljCdTUiLjMo2Mb3R94LkNqkgCFYtkgbFTmle7BrmE0+ZaxqVoIRD1wZSHZAQxcuu10512NJIFDw8PmbyRLOqKhZVw6nUgR85B65hqiQPRjn5fEXwYYVAwp5NRuEv9nFNWqZhGsNivqTIJDIXrDUsNjWgUcpyNa+YPN9R7YKQvXxRMV80zFcW4w0XlyUiWaO1ZrPZcnlVslx7stpxeVmRpBuSRGOM5/Kq5npp2a4s1sGucTy/WnG5MWysDF6sFn9FDDAE26CoLg4qeCkFvY8x0G2gdesMprS4QR0t5z2uJZUW4nvoCWGYn8T+GugWeKsY7MuOfiuKAyaw91Bf9sM3ov2eFYDXOxxEmyceF2lbhEL6kIHZplt9ndaLt/5M0XOy7qg+3vW/r3V3OhTqr+j4De0R9pXHgx9vPf7rtG6/K7xEBIyRnlAS1oFuDKoyyG2NWleITYXdldjdlqYqsc7ivUNqTVrkAbRoPEJMRqjJCFlkqERhlcfK6GbGI73Frje4+Qo2Jdp7ZgLeHY2YpZrW3Y4QeK1ZlCXldsu5ljwcZ6Syhj3wlptuz76Erg8TLzVOKB5tap7WjoWQVFKG41pglOGEMPwctP18NCIrcpTSew+z9aK21G1rS71Yka9XvKsF/+j8lKNCoSiDAuDj/r8P6aJOpTyrHP/28yd8Unqeq4SmyEhnOflIgzQ3+tSqrGkquXv/hB//kz/lw++8x3iUEpD76f1QkRjDjOx7LrxoI8ZVUIZeRVQ3aHCwnkQfsKqUYjQaBUVAasrdjsb1sLiJVp2Sud266GaOYkoSrD0pIdHYLGXd5Dy1nr96seLjLOXtu1NSnQWAoNa69i7EhNiS751O+PZqzU+XJZvVGrPekKYKIXWvM3bPFoSSpEXOZDKh2SywcespCOuDiMswWFolwANGOWpnuGpq5k3DxkpqKcmcwDcGYSNyouj302/OaetpsCgc5+OEiVQsNzuuypr3RIKQGhGhsceJ5nyUkAmL9hbpbNzCiEJUxDVNzO7ADISfpKkqnj96gt1tGBcJ85Hm4lnGOFMoLF8+3nDnzqOw1YVnuZjz4tkztusNSZbz5dMt0+kEpRVVVTOfL3j2+Bk6VXz5eMNsNkPpkP307Okz5hdrqspirWdX1VyvK0orYwpjC82+b5iE+JQ+HFyIfiN4PxkxxGQ472kaQ9PUET08en2to6kbbkZp76/2YZZg/9AFYfshxFb0JBCQEtrN0/0Uwb0LfKM1gD+QB+BVc3IbB4rBIV2o/O8g+npQ6/Bx4BIcktO+9f/1256FfvD5ZVd82fc3PQIvP+ZlHq6XtqGhi0c4F6vzga4Nalvhrlfsnl+ye/Kc3RePsVdL2O7wZYmr61CkR3jQGpFlyCJHTsakD+4xfvct8gd3Sc/vIMYFNk2wOmySSOsp5wua+RpZNiTOkzvLWaIZSUKAnLN4ofDOs64rmrrmPBtzlisSO3Rntlp5+3yHAVvQOaBF2KN8vFjwvHZsRLDSQunWw1QtATLWT4/oZ0LAdDYjz/OQG3+4zqOFILykWm1hs+PI1Lw/0nz/zpRCWIRt0/6iUqIk6IS1l3y6qfir6xVPGLNOcxgXZNMMtAtxKSJeP/BEHB6lBXfv3uH7P/geH333fUbjHKUG3hy/7+3ppqnjqOwTmb/lbWf07FOWGP7YXTv6kLzvvAEtR/XbHcaY7iytJd4nGNOwq+3AOg3r2wuBSBK8dZSp4dJ4PqlKfjLf8rDI+O75NHiJXBOXsA9xI82Wd8cpH01HPNw2rMuK7dU1ejJGJclef7ugyJjieHJ6xPpqiTWD+JG9AlCD0Q94h0VQK82qqrlqLEvnqaWmQaGx0LiAe52qlyzQobfGonzDLFHckTmP3Ia5aTBIlIj1BZylUJo7ecJMeApvWWMwUUDt3yIoBFILRBKQRj2AA1sZrl/MWWqPkp5Ego4GVpo/Is3CVo10UDc76qrCOoOQkvSnX5AkKUIonHPUdUOzK8NzL74KcR5x7dRlSVN5rAseWGMtjQOLxns98IoMCTPO+GCZv5ZP+qAEtABYrfXuI016165ph0wEKlEDPh//uhAQTotCGGnLR1roFKtu7fR9HToJYnfiUv/mAgT8nhWA1pp62Xy0s9eDt/QOofb3ry+Y27O6QI026njvtv7g4fn9n/8A7U2VkDag6aV4OLc0Pwhakd6jrSetLOm2xjy9ZPXoGZvfPqL68iuai2vqi0vUpgxeAdOgTAPe4qTASUWjNDZJ8GmCPjpid+8u2YO7ZO9/m+NvPSS/fwd/NMGnmqRxrK6WmOUKWdWkxpF7uJNqRtIHpo4HCTWOpWlovOW+UhQKpB2gqw2BXobWlA+WDh39SJwXPFnvuDCejUwxUoPvQsQPJ6hjYAgQSjGZToJQE33ecLhtyzwEzlqWl9eIzZp7OD7ME94tNKmPcL8OWhe0J8HJnGdbx3+72vAbI7lKFabIUJMRukg7xMeujG/L5IXj+GjG+x+8y/c+/oCj4zFKuUPj9uawBuProLkirceqwf2xLQ/l662B1huglCLNAAo8jt3WhXQs2uwARVJA7Ry+Ae9dNz6PD1sBOsHnBeva88zU/HxZ8f6o5IPzOyg0IRCtVdQcNDWjLOO9yYj3FyVPNhWbizn5vXvoUYFEdBzIiUAdUoBKJLPjCTpVUDbsxezsAUIxUFbChHkBjVBsEVzVhuvasis0IxENF2PDK21prU39PHhI3gfhJBxSOk6yhC8ULKxlbRyZbFMBLVp6xoniPFVMjWWOpRwaL52XwiOUIC0yRrMxde1oKhOC/1xIVW2q4CVo00JBIGTV6mIdCFFrKoEFYSJOSvCQeAfCxUJY0oTCWG2WgXMxc0LSxveH6n8G791AufQ96JDnwB8rursPCG2fbbeCuvX6tcd0/D16R5QkG2cU4yyEkXSOgdsovVcCWgroJFirjItB6MHhuvtmhwD83hSAlkPSWlUvr5Mg+jkXkXkfuGq+douqZEvgr7zOLRvrnq+/7QC/uxfh698o/Nkz5oYKzC1YBO04AyiPJ9k1iIs168+/Yvuz37L69ZeUnz1CP3tBXlYcmZqJF4wl5ILIRh1GSCosG1tRCkHloHmypPr8BbvZl8hPHmM+fJfZ995n9ME7FPfvkDvP9XyJWW+RjSXxnkIIjrOEXBL3/z1eStbGce0sRgqmqUKJNljqEL996As5oJa4OBvjeF7WzJ1gJ2L636HK3p2zfx2VpuSjAtVaNr3PqD/VeZpdxfryktl2xYNU8J1pxkw6aGJVw85M0CBSrE/4arXjb642PJUFqyRFjkekowKhFH6wl98GdgkBSSJ5792HfOc73+Le/VO0bhW64XgG07Mnw/q5Eu04Bgphn90xOPENjZhW+Lc0F5SAlDbWpixLrA2VBqWUJKkkbQze27CdP5hzT1C8ZJLSJIZFnfLbuuSXq4o/3Rju6wSFgpiHHmSTRXjPw9GI74x2/HS+ZHm1pNlUuClIHQWwCGP2ERJcKEExzkhHKWJT4ZteGQkHDDWjwZvIqwySCsl12XBRNVSTDCMisqO1eNOCLrWLtVWt/P7z6URMzazQCK1YWMN1VXKSCxQevEXgyLXmXpYwNYbUK2QrjDtvZxTmSpAUGaf3zwDFarGlqZooyeLmi4+YEHKAp9HJTk9XkKkVzp1NJjs9XPigADghOoVMtHOnwloTEJQEhkk8vVLrBgr9Yex8q7S1HjRxcFy7PoLsGJwoAOHw0iGkZDQtOD47ZnI0Rsh+MIIBrxw+Y1yHRhu4Xvgb1LE+duZ3lk9/wPYH3AK4bboGi8HvK+EtOtf+Ht6b3Sq4+9tkFtm7KtmjnH+YTxDamh6vnBZ/y3vpPKlxpNsani9Y//ILnvzlf6H52W9Rz68Yr9fcqUruO8d9KbiXKE4SzTRRKB24g/GCReN5XhoWjWXh4NrUXNSWq01IhXvx1WMWjx9zdvV9Hv7oY8ZHRzBf4coqQiJ7Cik5yhIyKWjBcbzUzCvLtXM4rZhkKfhWkA4tqOHfg7QtAcRyyZuq5rKxLEmppArpf28wW0IK8lFOlg/y6feOjZjpxtKsN5j1isSUPJjmvDPLgNb69/R7wRpUyqa2PNrs+PWu5iqZ0GQ5o6JApXrgmGiZeVQ5hODkeMaHH33Au+88IM3U69TawajC2hOA2zNP9kFew1dD8JjfrQVoYEWe551ysN2VwdoXoKQkzRKcd3hvArSwaPfMg+EotYRUs20ynpSGX+4afnq55PzhBGU0EPd3W0vBee5mOd8eZZy6hq+2O+rVDnNiIjxw7FtnPXqElOhEU4xzVvMNTdP5CejmX9DmEh9MrMDEYMBFXTOvGyqhI6StDMW+THz+6ka8PjeUtjbQL0tQWrFuGubbLX40iuaqAWHRWnMn04zXOxJnkD5scQRWF7xe7UB1KrlzfodU5+SjJdvNlhYQpUuHFiKWsh5I+BgX5JyNEOQy1CsZGGadR8T6mGJKL1S75djTbgvbEZTCoSot9mDOZUee7VMKmS89be0fN6ReJ4brhSDApUXphJM7xxyfzMjHBe0Wwc1nGv8THlQ41+IiSFLst7jFc/gPrH3DsgCgTWtq/U+tnieECMFabzjnQ+1QeRG1RBEv2/7q8NLuqZo3UEOHF/uGtjdz0Q4RwsIiTK0j31aYRy+Y/82veP4Xf4P/1Rdk10vOyor3TMVHyvLH0xEfHY15Z5RzmilGWsSoZo3xMN8ZPl/suLSe543l87LmN7uaz6s1T5uKed1Qb0teXM5xFxccff9j7FfP8Ost0ltSAXmiyFOFViKk95CCzFhWDWvjGKUpp6NR8A60QVV7W0MtpzkQWDEAsPKSrxYbrqxng6Ju08j2JvI2Hx4oLSgmGTrpA8LEwRaAB2xTU66WZE3DKfBWnnCvSENwmrP71xYKpzI+vVrzy9WOF0Kx1glqkiNzBYoO3nX/SXu0Vnz4wfu8+/ZDppOCUCClXRjtX9d9Gor5YLkMvAqt6iAcVvQzF8TH351GLKWkKAqstRjn2O1qYn4PSZJgvaPxFiqCBItBeF4KrAZyTd0kXNUpn1YNP3m+4F8+PAoBhU7Rm30SrOMoFbybpbyf5nxqbIg5OTuhmKShHHE0Y3urMSgBxWREmi1ptluGVvRwVjo6i9Zv+ElglWJrYGE9GwsNIY9eew/W4a1BaNUrpnuz3ZrbMjwkYzktMqaJ5qJpWGx2+PNpPC4EpSbCcyfLKOQa3aZZeIH3EuEUsi0SFXmeziSzsxnjozHWmDhnsc5K7IpqlVkpujgpicC7JljnQvaZVTIE+bno2eq2EERUMaPC1IlvMUCe7GY9tuiB2LPcO/KXg69cr3jsPR3ReXNalbyN7xeDuwmtSBId9v9lDzYcIINFlPcyZot4SER4SaKmEdPRI2z7N3h7/43aN04B6BbGgUTr7ZPho/8al4xXOdxXEj3FxK+GaX/i4Pz+Oi+7w++7vfGdB1q49h7tPPnO0HzxjOv/8guu//K/wi8+4+RyycN6x0da8qenI/70eMxH44JZIiiEJ8WgsGERigRvPaOmYWQbVjphnma8V2R8a2z5dVnyybrm87LkaWNYm4Z5veVvn10w//IpZrkmM47UeUapQitNt0MrFV4lrJstjbXkiWY2yoN1NNzSuGGhtky6jyMJ5X8lz7YVGy+D9S8PAvlubJP0rEVqRTEpEGrgHh3MfVtrwtYN5WLJxFreKQoejMYUiYS6hfxtj1cgEoxXfLna8eW2YS1TmkRSTHJUpqJSGjMhuuhlj9aSk9MZ3/no/R6OGDq3fZcC1nYwGnNDkhaH0wUxvjYy6dYKlK9A6/oabbgFlec5jbE0xtM0IVsBFazvxOoATmPa/rcmnoBE0SSKTZJwUXk+LxuWpSFNE7SyYCpoBZkzKG+4kyV8fHLMf3qxYrVeYaod+GlnVIR4gBb/woGQjEYFaZayYUu/VdBOnAyKr40O4EEgqhcCKxRbIVh52HiPiwl6jmCACGMhjwGng/XYCf/hc3GWaZIyUSkXux3bqg737B6mI5Geu+OCqYKscWjn8MZgSgOjDFpx69s4IR+C33Qb+0JQALqUWrpMkb4AWxSmTgU2KWRUoELZcgt4F3AWJDIORfT1UHwvgNtHKnwLRNXDoouh1yGe6OOWQpgqwZAYh2y7M+fa7QwRgeN8u+0bhX8bG9HGBRzKmKjMGGPCdSSQa8QoQyStN6XNohHdsxARfOkfoi7w96oAvE0ofGO+Lh8JKln3MbxrMz9dIJ6XwD++vt0mLET3Maz1oEnLV95hIGC+AS6Cwz3/YVrWcE9XeUgsZJXBP7vk6j//nMVf/ReZpH4AACAASURBVBT3t59ycnnNB03Nn+WSPz8q+OHJhHcmBcfSI7uI6ya4IJEILOwsadlwbD25hInwnEjNeaF5Kx3xjk742WrHL+qaz1c1V19UPJ+vabY1clOTWEGOZKYVSkbBHRmuR7AtK0xjydKEUZJ2+AC9GXGoELaf20heiReKxkkuy5rSC4ySOCmikB1of3sWugx0IBUq0YxGI6RUNxWOyMitczRVRbVccW4q3pkVnI8KlIgCY8jgpMQpzbz2PCprnhpDlRSITJPmCUoxSM8L1/eR6WdZwbfee4sHD8/JR0kU2oNuR0XDd4y4pYluVnpjc3h94DBH+ndtw2yAw6a1Js9zqsZizLYDn5JKoZMEUceiNy2LbwWeVpAoqkQzN5bntuaz+Ybx2ZiptCBauvTRS9RwlMB3jkZML65gt8GWW7w1oDXtHvLQ6SMQFEVBkqZB6bBhzttf96X0MAc8KAdGCCoUGy9YW4+TKmSyyBDzgGlT8rppj+d79mICvANrSXVCrhKk3VGVdbSqI79ynkQJzsY5R0qQN8HTUDWGzWrNaJqRJBEdr+OnPZ8LNBAZ8+G2xt7+fTxL9vx2KEPbaRLDa3e3aG3/ofLb/rZPGxGvj6EN3xfmvEGwHTphf0vRBbMKIVCRt+9jXbR965WTYcecc9RVzXazC/3QEj3OSY9GyDSJ2wqht8MOBaC6NnzyH1b7xnkAggETrZ6OCVra8IveF/Bq8fyaO8R3BwqAZ2AevSkj9Lce/XdGCLd14+tcvPexdRj8WWPR12te/OQTrv/qv+H/9lOOL65531T8s0nCvzmd8oOjnHuZIqGKAWyerra5cOAicldZh0h+AnxvYi2FbJgqxR2puTtNOZGSyWZLUlX8arNjUTYIp1AWUgsjCad5jpbyRufLsgRjSWWOVirA6Lo2A+BAcN8WdNkyZye42NWUXofCP5KO0d2eBUBgthJkkpDnOUreRnPB6nTGUpclZr1mbHa8VUy5k6dxP3do6QkQCoPiq23FF1XDFR6TSrJxgU4VUraZ/PscyntDMUr44MNvMTsq0LEi4EuxH/cspnCt2xLFuvG2euKeInTz0Ne1Q8E/VEaFCC7/YpRTNzV1Y7rvlQrKljX2Jt1LQGuMNmyV5EXj+enzK751NGaSRZCc9r5RAZiohHfGKRPhUE2JLUts3YT4itv6LSBJk6CISIW3rp+DvXnwh1+AByMEtdBsrWRpLGRJUACExGFRxoBL6FNWW4Wi3dKKF3IOhEWojEQkeCvY1UHp7qF+IRGC0yJjIiEl7NU3TcPFxQuKScb/z96bPkmSWweevwf4ERF519EH2WyRlMTljMSdoVYyzdqu2e63Nds/fGZtxrQajUbiiGSzeTXJuiuviHB3AG8/AHCHR0ZmZR/VLFKLtuiM8nCHAw/Au49Du8I2ElNdFCogTf4zkwNoxreJ4mqYMdeaTCUTicvjThKwzgWnrOjP13b5QJ04rtTVDkswMveyF9TTTbm/zAJEpl2SAJFneeOxpOrX4ndVpd/2XF1ecXl1hdcAldIcL1mcnSBNnYZTbob0BpUvngL+99zeOgOgI9Z7842xSYGMlIn4F23nlvsDvggpHM+bjv8cN/IXbLu6hXeqafQgbgO0647+l0/43X/6e/Qnv+LkxWs+Hjr+dlHxf334kL85XXFqXCxXO6R69SarPLNYYGIiliHa5I2tqFUx4qgCNMHQiqNpGtqjJW1dwcUVw9U1v3SO8+Tf0WrgEHi8XNDY8h2g3uO2W2oXWJjkFFcW0QHmUtku1HVk6FxQnm96ulDHbJC3IpbpURTEGExd0TQNOaNkVgOORE0V3w+4zQa2aw605/224rSuIGxSh5nRiMmHnBp+cXHFZ33gwlpCW7M6WMUkQ2aCwdRisZ/Dg5pvffw+TROjEWRESgY0vGH/3jbphEDLKmtvMYLFWkPb1izbljAMDOncGRGaumbYDqjuGasVQmXpreVlp/zTy2f8H+5D3lvapIbV6RMcbVXxYNlyYisa7wldh+t7jC5ubhlJWpOqom5qbG1xPjDliLgLsvGdHonhgEG4HgJ6sEAxBDGxkI/X+JnlkfAF8S/60xDDIG2FAzbBTcQnma+sBI5ay1JIiYfBD4FXz1+yXC5QzlgdLbB1TPsc90oYGYDRCVQn4ivZJpri6VVArEaNq5aZBuPf6BCnU+RHZiCyr4RE7Vd2nI3KjgRPE5kLyQwIRAdQpnvLJZpDyE64fJehSBqzrCXQlF1Q1YAJk0lNExRU8W7g8vUlr56/YrvZxpc3lvbsmOWjM7Sp0JxDIUch7NFw/aG1d0sDMHKZBVGeKPWcE08M/+ch/jdJ9CT5S5j0AV94+PlgvIV9UaK3N47jBssdlWGVh7rz+N+95Py//jP86Ke0L1/zQTfw123N//3+Cf/h7IgVQ7RbuyT55+IcACSHKyq0HyJCS+lGw+hXb6gSl3Y4OKqwxTY1cnwICvbikk8ROjUs1HNshdNlRWV09ExGFYYBHTasUA6M3QFsyYxQSC5z6TV7jgxeuXQDPZoQgJno4V6gRiRoTEXbtlRVdQsbG18evMdteuzgOMbzqKk4rAz0KVVtuVNFcCr84nLD75xyZRt8XdG2dlSJ57SoeYCK5+iw5cMPHse89SkKY9Jh3SPgOPUtNwhOoRnQnQJAb6EJUIvhYLlg2GzxbiCEgAFqW1GZCpdr2pdhWdZASjF9aeDTcM1LHfgYS1sSVLFk9G9szWnV0HaO7WbLsO1pApEo7IlwMMbQtA1NU+O2/SStl1EG4ywong8EUXqEa4WrQfGmIkhKLIONSaAcY0jc2M8oyeg4btSAUUxdM1SWCxJTNJa4BkSxVoiKs4mYM8CT3zxhs9lwfHJAu2yxUs+YOhn/X9jhR3hManNJaxDnMD2nTPb5WGjplmDp1KWKHzUEoiYS+rS/hXSNaU/DhPtL88JkVphmEM9xmdQ6agNyNEP2HRtpS2IWNYWBeu+5urri4vycq/NLgirUFnn/IYvvfov2ow9wTT0xYAriNVa4/Fw06N1r7xYDAGkxp80WEy7KhNwLweBNQlzZpeaDo4lASrnFJTq3kLfJF6TgaUBvgy/cRTdzIv9mKNgAlQ/I5TVXn37Gs3/4F6oXl3ywXvODxvK/Pzzirx8ccaAdJhP/3VzXmf1XExFZ7+KSGIMaKbQp8RRXEitlNX5AgL5u6E6O2HjH6/XAa/UsCBxiOLYGO5p5JIkXHotjVRmWdZ2QSbYP53HdBu1IwLNTdReUDTLZ8eKmYD9Vz9ejx33bLrDWpphhijXO2EoJg0f7nkUQjqzh0Bii39AOQ5Jg5Zzn6bbnXA29raGqsXU1FiPMQ5tCVT0PHpzyne/+CW1TY8wkJUnR/53tzo1piNJoPHHjI4Xq/r5t371z4hOT04S6pmkaBudw8SbqVF3Q+yGGCo6nPEm+1hKsZWuFV0542vdch4bWmmIt09qjGCs8XrYcdD3rzZZhs01FqsxeeBkjtG1L29Ss1YNUjOucowx255fgGoBe4Erhwnt6wItEj/pAfOeg0NbEA1QmBNqVHmKZ63q5QJuaa93EyoLpDMaYe2gtLI2h0hxlEvvzvefi5WvWFxdYaxAzZbvMWiwSXp2k/2leZWhesYqzX2VU+afZ39hf870/Ph4kbdyQOYwIm5EBKIUznbqSckRmZ4xh9sZJkNy9L889MdmJCXBDz+BctP0vK+RkwdFffo+D7/8Z5uEpW5tY7FHqTIdUJe3TfS2+15h3txrgW2UAQgiSkvh/nhZ9l3R+AUpkGP/c1e1IKIWxyJQmOWlPSmhUJN1X/jjddROp7UFy80e+njaTSHQ8QHOIKRXQDo7h6XMufvIJw88/49F1x/eC5z8cHvJXZ8c8qAT6bXLCyhx6ISaXpTn7mN1MiUQtjGOYkIQIxCKfgYUqDzB81FR8d7XknzeOTfC04liI4bCCSnKiqHS4XEA00FpDW1mmsKviEO622aU4+16V6+DpELyYItuYmTZDiRTzsxKz1TVNgzGG7CQ3amJEk7Ze8UOP23YcAQ9tw1IEm+3/4zsiEfMI1/3AeQhcYwhVjakbjK1QSZ7xwmwcxloePDzjw298gGSbbh7unj23u18jo7BjZ70BOLntx6+0ZWc2a2NUQC4YRPIOr6oakZIBzbXuBaxBK4sTQ0/Ls3XP9bHnQW0mWGiSpFWpBD48OuH0csPzrmfYdmiIDMiUZX4Oh7quqes6WW0yIcpSu7kV5gFhMIY1nnM3sEVjaGVeUAVcmPq5E85xrzRNQ93UbLtrnBvQ7EJAVGtXBg5tRUvAhLQzE1fonce74ebSml1mKf8mxZBuG5tO9+KZdJP7iOCbhJSSezXFfcW9Wegrx3ijv4kBuNn2MTDF+7PJ0QRoLLJcYB6csvzexzz4D/+e+jvfpD9Y4EyOZYj7dHJ0zePNmpl3ltbvbV+PBuAriCYqFFLx2z1VL1nbG3Imp6y2GvdRFLWmPZZJ59RmhH0kPDsI9saVr7bduq32IqNJHZdRXB0C9abj8le/4fKTn1O/vuC9vuffrVr+6mTFx6sa/Bpc8qQeiX8+WGlzZ9zaO1IlTOaW50k9OR7woFgVFjpwBJzVlpVArQGLp5HAqgaT1YIZkINHVamsobbF+0e8rcxj3PY1wxDgygW2SMo0Vhzavc/K+KlMRVNF7YMm7j8OIbFWKcbb9w7telYivL88YFVV0XciFFJeYgAGFV53PZchsFVLsBVV00QGp4zR18w3eJq25uT0lOOz0/h2zSGt99t1mSm8C1XCPkb3LbQ0LyORwFVVFbMDhmiPrasqOkLuG2jWAohFzYpXmyGWy21Kwpw2afBYVT48POTM1tg+MmlBy1JRN/dBVVVUO3UDJiRf/DO/KjkgBjEMYliHgYvBs1XFFQIIEJMC7douR5iHGb8NQlM31HVN2ELXD6xqkwTYUZzhoK5YyIDJCXkMsKzTcNO78rlKzpRS19Nv5XyKC7uWonjktPzHCALy2b0huGUGSilNpNENQO58/9h5wQBk6TC+/gvu1QJnxuVTWNRUh0vaR2csP/4mRz/4Hqv/6Tu4B4dsqxjKeXeHO0zL+NO77SjwNZkAPv9CzaE2P3wpyvNzDiEStWhvut+Q7o9e337b3UUTB3rzjkygMgtgFCqvyPWG7a9+x/ZXv+O4H3gcHH/18Iw/PVpwwBA97MeEOpn4l1g4nRyv0A/J9mdmcJrxSTqNwapSozTEeuZWPUI0EVRiWFgTGYCR+SCmUAWMNVgjsyR/92sxFeugwpWDLYKSVdx7VnYkHhnG0SZc23nCINm5NYSADh7rAisRHh+uWFR2umEWf2zog/By27EOSi+CVhZT5xDDaShavKdtWw4Pj1gtl+wC4j42+/uATXbeP46dt3AOEoGrqoq6rhmG6AdgUWpjqazFBb83ogCJznbBLjgfAlsXiNXaSm44kCvrPWxqjo1S9QNd36dyvzDmi9A5NjHWJGfMYk1uA2COPkiRJQHofGDjHT0BZ8BrND2pgKRCVxi5VZMwQjtAYy11FUv9dv2AP1jETHwF8VtWhoVNGicTwBoW750iqyaa5rILjwDWYA+WVIeHUQF2I7lasQd2hB0ZJWamM5pZ4cxkFCrymIMgdZ4ZABEkpJz/JSMkM8yRV6L4rgk1CGqSp78Wa3Njg96xYwtkpUaQymAOV7QPzzj68BFHH32D6vFDNquabSXRPEVKFJTP8ay7mYqiGHFKL/QOZwt6+wzAPG7ino8Uf2+I34YvzPmlriRpfG7tpTzzymwCv6+VvPO9eyZSRi8bVYwL+PMN4cUl9eWGowDvG+E7B0seNAJ+E52Uxid33pgl+qBTcZPbcsWNRGNS2eeimWCi1y353CoWjxWP7B6iFO5nJdpmx9/utfx5EQUXhI0XOmq8JhOGlgS3QGwlwRmF9p3VnyGciMjEO6rgaIHjxtKIzsP/8kNicApXzuPU4sUQrCCVzPL+z94h0LYNi7ahSiVlM4RL4m+KR/ety+61fXH6ca2SZFcqc77illn4XDWw67opAQukiAsTi9bEByAln8EagoFODOf9wNZ5IirLcE4fjSako7piJZ46OPrgUHVAPXa7S4eNMRhb7o/7obBcwjYQCwB26pMGQMePJRAzHSYmVHffXrTgqalYiGBQhn5AdcmYiyLEOS6N0piA0RBtQw28/71vU713ylALIR3DYATqmoNHDzn64DFhUeMs6GgS0NGNQEjsvwhGcnqgsCPQploKks1iMZYfmSsfprsjE2Q0xnbt5p0QySWAJUEzM965XkHMw5R1ajncb3rLDOvdsWKTGS8yABZT15hFA4sG39YMdU1nhSBhnEc8eXMtkEgWWEL0BdhNaKT/in0AYrOfi/rvEn9lX/ptmd07v7qnQyUiaSE6ct2hAx3lh/LsF5q5r73NXrpnxjPNk85uGcN1AHxg8/Kc/uU59brj1Dm+uWh50Bpa8RB60FSFb5SQb75PQ4ihgTD6U0zvk0nS0PlzgmA02t+jaTx6/RoUK4oZY/LDpLvw+TyZuIvmqrVbAFUS6wgfp8omKD0m+gDcuPcW+6VEhBoJoR+tDTuKAsQr4gPWBxYox1VFLczHG7EFisUFuOg9TlLGNCNgBS/5HaV0H6G3XC5YLJoiO9/tcv9dQuXNe/POLiQ7yR7ltz/35drUac4LUFUVXdclSdFjTCImM3V58g8Rg8eyxvK67+myXV2i5zyj82D0PzmqhaXRmCnPh6ixKaCsxf8RTQxAomKaz8M95iORyHkMA+CcxiBmyWaAxGhqigqZCTe7Ld5XiaU2IKoMziebcyoLrAp4GgutaAwFFMAK9dGK6uwQ3wrepsEZgzOG7mTB8r1j6kenDIYxxW98a84EyZhCOCOSnLlPNF4PiejpSOlz7H/SCiYNYSbZmvuIyYVTzYcSjIkJGWGaHbN1dLQbTbg6nYNpfSan0VQ26ZYWxrkoBq3S2RSJTro2amwiNkpvGdFJdoBM5y9HbmjBzKSwyAiKd1f6h3cpDwCQbfFz1RAjo7xXXknXd30Cxsc14oRY6lRvU/7OHlJkJhxm/PhurORuZrL5ldgymZomIcGzvrigv15TuYETdXzr6IhVI9hUYzx2UnLUxffEROEC6oYo6Yz3FktcIgtCkglibm1BkGBSWvwoiYsYagINBiNumoEqznm8EuOhd5MEZSo8nq9c17NcpXgoB2AdlC0xWUtEeLJf/JsRmxATAtrd8r/TGCLfouADNgQalNUuA6BMRBWJGoC+Z1AlWBMr3qXY7pCRaUa+GvmDVbugbZvUWWC2i9PX8Dk3aHmmZI9TzV1x2F+m7TI5trLYKs4/g8xagxGDzyGUOWTMKGKVYGFj4Dx4tqmwEKOZKIeDxtK6K2tYSjRDqdfompFhkCY6pozVEEvZZgYg+cPeCxCancBs/KikkEvJDuOxL+/T78X+nVXwm5o1U4Ge3rnoUmKLUEB1VEaoRZLDbXLNqwzUFaEGZzX5QglOlI0MVGHL4dIyVDWeKUJgjkSzs9u0VtlnLjsijvn3I1eQHjeJLGdYRG1hzvIXJfvktV+c15GpgOL5+MTkgT+Hz8QECKKTpf6uvHxZ/o8EPu27sseEG8ocgjriOB3nHnFE+n7jValeQtRkjXLDu9beOgNQ2ejM/cYbR1tbXOQpjW3cJHcHWtwC3Uz0RwYgMQS8mQm44SX7ViShe7SdiU0S91yOvSEPC+OBEALqBzbXVwzdhsPgOJLA+4cLGgMxhWoRfncDmAJio+10cOAc3tSTd3OC6MQr6YwYT0cxHetRdWAwKjRiaY0plHaaeA1P0GQvHNWUuwd7Z7A766QCjsA2xLCsqJIt+9E9z2YsRxQq9/h+SQZLIGpFvMeEgAXayiazQdG35ggHxauy8Y6BjIAiAxBKYJXSkApt09Akx63x5935foE9OtVUmmds29f9V9YKnhLAWMFYg7GGEGIuCWPM3jlG87eiFWwH5cp7Bk1S2ZhHIocMR1txY4SaEElQCPiQCYuOmj5bYhKrMZXADYZyZJf2z2c8D+mjmfll8qnVPMZ8MSXNEbihaUj7DxMl8m5wcRvZ8gwolTFYSUVq0ngDkamL2geNZgDxBIQwdKzX1yzUE6TG5zOR06snFCCJCRVkcsZPjn6Z0GMMoz6luF+gEMoidHMIrklaDE3jLdFr1pSIaC5uHMdcnvsR/DLS3ziawk/sDnKbo4CiA3OBncb08nGOZTn6kOGRV3dkYqe9UO7XqKgSNVb0X7kJ4KtptyGi7Hh62+8lZzceGblhbf4DalP40rgZtfgtn5GkIjPJW1z9gLve4LcdlXqWohy3TVQb7qarhQnxSST+UINzaA/qLaGSSQ1WroCSbHlKdMIri2RkhDc1g1ARy8JKcbDz3bOZlmFKb+TgJik5aGDwYZQkZmaKGTXNcw7j3MVIVAfvfVMcjwaNaWNDhHllbHLUSuMZsVT8KOBQHDH0NEsK4/B3mRiNaukq26XNJEF/FUl79p6fr4npjSASTNKCSIL9mI1g5KMiPLNy0AODITrahRwVQXngR5DbEUoexU/5BW5RTJq85p97/rrzmcBoVFP+AU3G9RCTc+xiImE6ewqSyu+qgnN+lF6nm2MKZSOm2Avx/OXeM5OTn/KDo99uURegArWgKQQzE+8gmpIlzYPbRsV7grdmM1bJ6zItWWYCyowOfjxu00MqOXLfkDUysY8smJT4gPna5XeMDIdMx+7WVdJZfyOzIjs3pn4yzriXQn/EL+8s3R/b12ACmGSML9PGNNXltZ2/dzxd8uXvpi7mDW0a91h0Mzadfr8VDqqoU1w/wOCwwVMDq6rBjF7Qk61ujmAMEUtUUfr3EExVjGGiFPMxyXjIcizBHHnlmRT3ZsPjDR1NQh+lw9QYQrRLLUs2nNiX5rShn3MbZhUeMRmV7pz+MvtZkN15pvfti6XKznWJyPmCvxnzUBSPZUlshIaCEPZEgszvu9cUuQkV4athLO7TVCDkHDAJ1lVmjEwZsimMYmjRIszndujp/uTsSemnrRODx/75jzZcLc6BFNj/FgQiEn0OKmJ46458Ob0phL1zKXqankp7MJ8jLX8XIbI3dpp1SngmWERs4pnjfLNLnfMB3zncxmGqgDU2ahl2IZHBmL+PJo2Jycn5JSbY7Z/R6E6x74fiwTF3lkw3RAbqJmNxO9Tubpng3+hih4OMmpvEEknYvXtsuvtFucXB9t1rf3AagLjIe4jOTpsLAlqo5zKh23Nj8e8vnA3wrbZpzjcZoX1ovLx78sgXiXZFmdWQL5DsjddKdGv2muqEFFSMzIxP7y9JPBKi0CM6Esep4lfxnDKx2Ts8Y/lTfKxkVoqbpPySsESaZ84oORHIHWS+dyPNYZGnqTr/WYxgxIySVnBR1TxL7ToCamJGo2QqieAwfZ+xewmpz6TWr2ZvxuFkc9vk96LF/99mm3bopE3Ke2l3T02jSoQnPVchUXNgTNIfp71eYGPdu47z/TV7U/Lp2HsWdN/3kgODXIGuTE470/LkYjtj8pjdjvMod/ZoTpO9c99U2CY1MznjFj588d4oY6POs766YrVaYmgig1GYXkvscRMAWoLv3qzi7n2377D9As4oTt7CO01RAW/qv+wzAyo9MyPet+OKyU1N80Oze8e+VSSEm27s70r7GhiA6v47pGhjsohyGTOg7yvlJCSSU6uOqCP3sZf436JK/JyS1VfdbhL8m7/NELfIaNMSQEyFWBtDqIgqVK9jQE3xKV5SICntovYATeFEM3vl/hFNWvCMDjXa9GcsgkTbnWZP5IkKjdI15QHbgxjH1xaQKDCYSNzoY++zfbQXlZDtyBp0h5svxpHmJ0aQ5LQG4EORGmmMbphgLBpz4VsFCUk1nOZ4Y5eZiGx7N9APw8zcI3lyX6KVc5uE0nle9bfRcoVAk5ditgzF+Rx/jHPVFGtuVKlVaRHqBNMbZiyhCFHL7y2J7s7ZyTeqTiFdwL5cAbe1bFfO2qCQU46PJjVTUOvdc5R+yNtSdVJNU+7dYqzoVD4jvReJ7xV00kGMIIlaJ+cd1+fntGcnSNsSPfcLb0fVmNtnljSlpMZfXkc0yztxg9m6pfeRLuz96SsZ126P8w5lIh+amb1J9xc/+fy/fSb6y7avIQ/ArQnX72zTZpcx7GSGrnfZ9tten2hLjjBQLZBbxi3lOuu9uv36muz/p9zye8YPk0MLqBqMsVRtg9QWLyk9rvN4rZkzACUSFcbk9INDU2KekpmaZ/uaHpU0loyESxklx/tm5fqkUZDpIRFMkYhl13xwr5bW1wC1THXdJlfm24h/mk9QNIQoEd7GcwAYQZIUqghOk5ZjNu8JiVojLIzFEpDsfxEikZGSAGQko8p6s2WT09iOtdkl0cq3sGO/pkMQ94mOn1G602K9lUk3nAmj9zQ+sCJG9IsCZfnece8Roy1UYj0QMYjY2QAyn6GkQkmaCdI9iVLR8rnIzmMT65t7s8w0brMzp3u+T6djdEvIDGwauPc+bp8ZodbZVs4tsz/qPdurC0LfUYUD1KTwWzGMxoAC2WYzxNtqd+7hgul9o9NXvu/Nb7znfG57WVy3yMcFVEpGoNT66f/vBChfAJ2MTk5KTi9ROJ1lgiO3IPEb70+en/PENbMYdm5f5neMJdjbRo4z01AyGojXxFra1QLb1AwirBVebTuGo3rysJ+BUojOfzaW/XXJic5Ep5+gt0dHTznndVyebMc2YrDGpgMfJRavis/hV0nCE9FYHx4o42rnXCBv4C0jsrBEibsmpoY1GUHOtADlDijyIAQdM8dNqHkCcORRJXpDi2XAsPEeF0JBtLSAr2JFWNUVtWyxGpCUWMmGaswmV+5/9YHNes12u5lLSqpfmvjvf/7r3e+qidEaie6Ux/ImPUzMUvA0qhxWJpaR3mUQk5SqGDZe6dUQpEJshVR21iXT0swYkns7cY2+Lao46QAAIABJREFUGDfvn0pI50HZ7OpeDHTfeyZGMEfT19ak0gR540VTggsepwGlSmPxqYebxGtM8uQ9w3pD2PbgHVKXmRT3r//s2N0NkbfSIgbPIYFfTZ/75qQyYf1R4LrznBV5CG6M692mHffTa32JZi3yxbDUxMWiMXRkrvL8fF3mTHQzVw4pHJBUZrxEzh/wbi/fvCnx6Jem9LGynDUsDhfUbc1g4FwDv7m6pA8+U+eiJ0OMq0/SStdF+z/Zglh6HO8OImkNsuZGBVFLdMYyiJEY950cvgJKp4Eu+KlEqARElKoy1CJTjvNSLMnEYBcAmseQCUhML9taqAhUqrNww9Ef5BZ7r/qAD34kEEFTKDcBR1L3S6xTP1jLRuG87+mVgrnQaWwhUEngqLG0QJWkWe3DLF27JXmOBxAf6DYd222H18B9omr/kNrIADg/v5a1QciuhhUTYKnKSV3HtMvZ30JglLJTNMr1oGzU4k00gZkcBlYonbTs3nuC9zuJFUzxuTEDJomPEWnEr+ls7ZHGb4FG0ZeMCmYkpk0WU94T3zBoqi2YkVZiwEfTZ8FvjPqIEKB3+E2PDB4J5Xv1hkSUS/7qvefx1bXZUHS+EuXniwzrxnzyAbyjw1FjNT5iELW348R3uL11BuD+bZeDnzyw869fevfJPdSlMh+J7nzeibY7qDtYc0XwBoIVFseH1EcrXNNwbi2fXa1ZO4cXA7ba0QIkWPsQ7f8aiX8mn0Zuqf9NlkxKjB0l+qz4t2byzA4oPYEhTHazMaFHRta7dvi7FqKUFNN9tRFWldDgY7rUkprsk/QSE6FETUeI2YhmmtcJywsYi9qawVrWKC+6nm0gMVAlExCQFIFxUjfUOdbZB7zzhYf1PAUJCK5zdNcdQ+eRHciXKvQRURf/zcCyD3y/580dQsD7lEo1Ne9crBBYDEwg5WcSKi+03nNS1bQmO0mWt0cIBeD1MHCpSp+SOhhrZssyjiP/VSVkJ8CS8sxfsCMipv9pLIBaiaGxdcp5x5j6ej6ZO5oUsAkxA2JbNZPj7si0W7qgOGX0d6CyKWNeDgecJjoOV8Gq4LcdYXCFX/Q9NsK+W+7CSffo7j6PSvnRnU9x7cvtZ7nxkVFFtG+05Tz2LOpXUAjvbba3ygB47zPFvicQskSmsytzFFBIb58ry+Ldu0Jz0gwmPmMciXzJPfWW2k3AyqRyHFuUIFxlaM5OqB8+YDg65GXV8MvtwK+vOy4dYGpm3tNZ2nYehpyMw0Y7avH++ZtGVz/Y/YyE18da9pLvFHySYjSLLEFBffKuj8MIGYMqxRhvjmC2hxICrwwsLdS4VHAo/777eHkhajFCCDjnIkOQtRqTbBejKYyBusY1NZcS+N16zcZ7YjGZbPNNjFFQahFOFy0LY2JGeq+xmmBOEFPAMUgAMXTdwOXrCy4vLsf3x32phPTfZGm+iaAyVGYaMGVkGPYkAnxrbZLuY/Pe45N/SR5rtGtnm77OxiteqQPUfuCsaVhYWzCduQcAg1fL023P66AMtoo5380U734DTpLG43y6HIhqmB3b7mxC00c0OnVahMbYGOkRtAg7S1J0Wr/563f2pIDTyACIQFvVKYlO/j0yn11QOo01uhCgbcDKhM9mXQpGYwRKBfiuwzs3xvXfJSCVxPaWO/iiu2hKl3yzRRDts9nvYr/PP4J9cyoZi31YbvckRaEgqw7S33eNWNzS3r4JADuW1C6blBtZi3MgeblLZj6l0tzlvu/ZsoPPnQwASe4q1GYl4b8tFfHvs8Uh7iD7YpATOVRcJZjTI8yHj/EPzriqKj4Lwj+/uubJ1hFMHQlWAVgNGpOFqBCIlfWiSj/+HaVL3VmXzDzMbLoxAsCLjtEd0UQheI0le4OWWEDJG8cHxXudc2Ryy1HfEQtEFWuUZaXUeMxoCHrTasb+vVeG3ieiFTdGqSEVQIzBNBUsGq5E+e12w9r7yCyZ0e1q/NQCZ4sFKzE0COICrneEQmsx7nkBFaF3npevz3n69HkKUJB0bnTv3nzjfs0w1pxEZ/p+Q9vyFjd+TPns8D7XXIsSuAspKWzB76tKpHI+0GigpufBouagjtXyGDUGmUE0eAxPrq957ZXQtNRtM7q8xHVUdou1DS7ghoKZkHsAIfdF1JNVCJVEM47VRBqEFMVwS4jh2Ca1gtOAS6mOm9qkseYNKGCErQ90IVYdjJxCM6avHPnlApHFuBvBKgzdFj/EGiCjr9Wec5VDh7+Muv3Lt31vTdf09jvu6q2cT6nMucla5NfcxqKk+2TqMV99l8MA3zoDoBa5ETWq+7dQJrRTCjAzHqlZzqzPA87ElU985N1cbnxzIq2lbfxrlJDu2ya0NJ/fmNITQKKfgzOCO1pgv/ke9Tfew1UVT43l/z2/5CcXG66CQJWYgDxnH9DeM+XBTh3eCxLze4KAs9BZYSOBIaUn9cbQY9hmBiA/J7FMbkAYnDJ4ZUpYdNv7C2oxAilQi7KqYrSzDcrN53f+nZkLNfhBGbqUg31MqRZTr4wI04CtK0zb0GF46Xuu1eGNJAfL/ApF1FFJ4KCtOLSwIGC8Jzgf/SwyoYO0/yKTFIzw4tU5v/zVr3EuzEzicW/O5Z+7SNatirP00G4s+Ntoo7kiKH0/4P2U1yE7hY4MQGb6FPAB4zyNBlrWPFrVrGpbMJsJMgYwFgf89vKScx+QxZJ6eZDyKsQJj3MtzrnrPX0f89d/PihE81UNLIwQdWq5BmbSzFkFSeoszeMtW7mOBudjFksRoaltwbxKOquG68GxDSGa8kwFiwViTXY9GPuVnbdYBNd1+KGPig7JHCdT7Y4yf8E95v+FucU3Prrvhvk1veWuLzqUOW4tWqYLIzoQ1MhMs/PVpL97++0d8gGIbTzCO/Sm8C27l3PueIQ0fmzQ5NQ3ZxXnh2KHT0nMSOZJ3rX13N2kgo5hbzAJ4hLAGaVf1Bx8/CFnf/4x/uyQV4uafxoc/+nimh9dd7iqQes2mgMCMe5/6KPUPntPjia+ixCXDBw4a9jUlgsxPBk6Njg8MR1up4a1j8xARmoxeL8GsfQu0OeKb3lB9r6zhIwfAVQjHFjLkiiNSa6oFiv9zLj2yScg3uNcYNsNeDcnsCXTjyimsdRtQzCGa5Rzr2w0aTFG7748LocxgbPWckig8g7jAup01K5MnVcxTaoxvDw/59Of/4qr6w1elZB8ZCwmynRSTbDbAx0DozSarxqJ9uqsEs5xMnmF3+a+V1Xc4Bm6AZeiTLIGwHs/WwewSDCIA+sDSw0c43m0NKxqBfVpoLl6T5TcA8qzbs0aRZZL6tUKNdX87CTNi4igQei3A8N2IGbALNS5b0A8oorVwMIKh01FI2CCZ8xDmV+aiUe+OHJkpSwa92XvlM5FJrxpqqkuhQgqlqCGy8GxCQEvArbCNKvofZ1wX6WSPHcm00f++N7huwGcjyXS36K25672ZfbaXemU9jXdp+kqf7+LgIsUnocxXbLaVHJ5N2lDvnfxuabztba3zwDoqMi8/ZZbrt2IlvnygxkZgL0ObJK4YCm+F69/ZxgAufmRpOmYtJXTaLNm3VmDfXDK6s+/Q/W9j9keLflt3fIPVx1/9+w1v147hnqFVi0aDPRRKo1h8GmzjxjiJgRLaSGveBBhayqupeJ5MHy67fnp63MufaAXoUfYYLj2SsgV/URADFLXiF3QBYk138VM+UyhwKgFUzdDqABKJcrSCMukS4pD3AViATNllCidD3TdwOBckohS0SKdhopAZSvqtsFbyxWGF/3AlXMFsk+irAZQT23h45NDHjXKImwRN9B3fUFkZHyB5BDWIKyvt/zmsye4QUcsFUeqTFLwfDrFpMbPhHDznBPrnR3f9jDIX6TtQ7TjKFTp+360/6tIlP6dEnZLG6rJ2auofOAgBD62Sx5aS3NDpW6jY6aAGwYuBk8nFmkbbFuTlQnlgIymDHkhMPSOwYXIHN5LpIwAM6o0GlhJ4Li2VEZjrgedGAAZ798LraK7aI7rBkffD4nJrGLBI4kMTtBA5wLbEHCJmRVjqNp6ygZ4Y+y5Rkj8ri4yAMH5MTrmC0nSe3DSV/bobUf1TfLHV9H2Dqo0SRdap31Pv40cHV9h+xo0ABVmdKPMiRMmbWq51cpDMrPFo+RUCvMUm/dtJbG637M5LPDrdI764i3v0CzFZnBPuzdgGIxBD5YsP/6Qsx/+BeGb7/Hi8JCfBsP/83LNf3x2wWeDZSMtIQjBKz55/o/SkmhMeiFFTXVh/B7/Hc0n3ggbY7m0Dc9Nw6d94L9drPlk63ktFZ2xbBEuA7zqPa7M96saPbabBVsR1uridZMI6g2Xtn2qOk0zV1ojnNQ1LYyVIW/CMHcxoUANHu8GvHPTXXsQTFVbmuUCFi0baXi+9Vx0iWmZ7fXIAFR4vn2y5MNWOQwdZtiy3WyiI2A5nmJ8IhXr9cBPf/pzNutudD6aIBFGaTanPp63iYErd0xZKVNGGHzxdqd0pSmcVAUXlK7rRgYgaKyU6AY3JgWaPoK6gLhA4z2nAj84e8xJbbGj70Ria4wB29Cp4XXfc+48g7WYtqVqKkZkQqHLSvP33jMMPS47AU6ZxCYENZ8Qeb9aVergWQFHlcVqmEJYi+QcYsyYB2M/tcpcvWXbDQx9H7MdNjUikw9LCErnHD0hVtpLGSnbZYtam5QNhlycK5/RuO6CDSBeCYNDnUvRN3NG8Q+h3XBu/ZLtfng/nqVgtESz835iX6LRB+CdJCNvPRGQJdeUmrDMPiJeMnaqMmn/AJJkK9lZ6QvAcnpb4nJvifuebtHfmzrs87XdvZXZ/vg3EqwUimSEoba0j844+8vvs/nNU9bXjt91jr9fX2OfXqLVkh+erHjkLQ1VqoSX8/VNEoqoTklJmHQrkcQJXoTewJVteE7FJ73nH663/NPllt9Qc2UqBGEbPOfB87Lr6UMbCXyhhm+WS4bqnG0YorNaJqg5n3qxR262zJ0Hamt51C5oA1iNZPNGhM6NLqJneRgGuu2Gg8N2rzQgxJr2zaKlPjhiu1nzZON4vR3QZbsjZWtiABzfOmj4uDacqefJ0HN1fY3rl1RVneBwc53X1z0/++SXfP/f/DmL5fssllOJ4Cl50N1yZtlj+ZKJRZ8HId6AzZdXC+A12v67riOkEFCviveBYRgSIzTBTbyiw0DtBpbBc2aVH7z/iINKIAwJtkk9JBZszbUXPrve8lrBNQ3LZUvVZA3AVB5qWh/o+56h79EU+RGRQA69m89hztgJNiQGQAyHlcWGMEnaI3OmjKqjzGCM+Qtyd9l5VBhSAa9la2I4yxDGPoIq636gC5pK+sapV8s2pQ2cnPp2C1mNzB+CDgOh7xIDYOfn6r5Luufa10LxvsBL7ox0+FxdThUX44PTk9nYMnN2fwfb288EaIEh046M1MqgjqQlKRB4DFWJquf4Y5Q2pTxAb2gTCczSaVzaKH1MfZQ0fwrV+WNqCQpJdHXGYA+WNH/yDR79r3/NkxeXXHcdv3ji8Nst68+e8Lp7wJ/VNY9lwXFtWGigUU+dwpEQSdXOIkSLAL9E+A1bsVyJ8EwqfrZV/ttlx3+/2vJzL7y2Nb01VCr0IlwFeL7d4vRwQo4oIoHFokVqQ++HKKU0NtUBkj1Efx9Tp6CBSgyPly3LLiYEmtiVgmEaN0BxTSEMPeurC07PDrAaCcgsjzkSExy1DcuTY9bnr/n1puP5ZoueLVLqWZ/VWaCKUc/jtuJPFi0fVlt+7h2vthv6TYc0FrHVjEnNR6TvB54+ecEnP/2Uk9MldXOKtRP5L4nZ3nOi+77m+Y9Tnsl/9z4Te268DdkG7+m2Hf3gpsc1eeD7HPOZ1jiAeg9uoHEDxzgeW/jO6SFLYia7SQNA1LrYiovtwE9fX3GulnBwgFktkboaM7VDgpcqWd242WwYui0ERzQlaBIv7S2AmF+sCSzFcFCZaPufIRaNkQpjzYtdxj1pMHIGTg9hGKi9ckRNjtTIONABrzvHOig9EUuKAbOoEGNSIqAoocbsnJlZz/+PmQXDMOD7aH76MuTqq+QR/yCa3p4sbtQgvOPZgd4yA/A+qoiRpGgLu77KO01JCrl4YKJ6MmWm1lIuuV/LDHbO9ndXy7nzx0RbfxQtSzBT8wa6yqDHK47+zZ/Sv7zgVVDWIfCLF+esN1tePTnnzxZLvn+44k9XDY8kOlytjKdGU5Y6E7PYkfwFRXAiDFRc2YqXKvxuUD7Z9vzjZc+Pu4HfasV5Y1kngoVXeoFOA6/WawbnoUoMgETpu60qrDH44Ol9z8I2pMxG3HehRAO1BB4tW9rXW4z6xEyON0xw2pW6A/jBs7la430Y55xbptEiYJua5uSQl5Xl11cbnqwben/Eom7A9Sm/QdKRhFg29uOjFX9y3vGPlz2193RXW6rFIvo/GmHMT08kptFu7vgfP/oxjz98yGLVcny0jALjDjg0E51xOnNT2GTCifUJ4jFLqZ4zPzA+Pqpa3gRtdqp27IxJISi+H+g32xS6H01MPngGP6RslsJkygowBKzzLIPjgSjfWjYcLhtsv02V+4qX2ApPzYv1hh+9POcVDeb4GLtaEqwQcgImZSykYzQCrLveMnRprbKPyQjcPUikiPA0KA3KgYXDukJ0bqLSrJEyWQOgRScZxgkLiYk5OEJPjXJg65TscGJSBzW82HScB+jSumENVdNAbVIZj2mDShZ+dt7mnCMMDvGKVMI99N/717bo94+/Zfdbzw192x8Q/fj6agHMz8+te6SUzrN9LlAmYPkC709OZW9K0PDHsXHnQZe79CxmBlT6ylAdr3j87/8tFcJTI3T/9BOePL/AbXpebHp+N3h+tdnycVvzQVvzsKo5sDE9b61p82jAi9KLsFW4DMKzreOzbccv1x0/6xy/0ponpuKytfhlTXV8QOi2hMs1Th2Dt2x9iAVNQs68FUOqjuuKlTW4YcvlZsPiqGXmmT0jTPtWUEEdDYb3VksOzJbWO6x6XBmOmh8taVeSokOA9XVH3w/UywqrUtyXpTIwlaE9PmCoa14h/Hrb89m6409PlpORUmMmP7zHuIFvHa747tGWB5cbXgyO66sN7mBJtWyw1uLxWBh1FhDH8/TpCz758c84PFiw+u5HmNamgINdqXJH2h1bmN9S7plStS3lhftitvl984qD0fFvs94wjNK/pGyAjsG5ZCkpQn5cgMGxGAZOXc+3FsJfPD6jUoeEAdSP/YCAsVx4+FXn+HTo2dglhycn1MsF43rNFjxlefTK+nrN0A3pJ2GsAiiwd3+N/s2KBKVV5dgajusK69cpBLmEZyTSI9OpRT/5neme0DucHzAWDpqWmX1eDENQnl2vufKBDnAGTG1plk3ymZwiK9B9dSOi46PzLjIBISTXm5wyPeWIuKcj2zsXUvYW25zJ3RFpJ/wh8G7nAfgaGAAd6f/9H0nnY08CDtnDTdxnBLmnr9JZ5N1su5De4cs17ssgMNSW+r1TDv/iTwk68NooVz/6GS+eXrBd91z6wLN1xyfdwPtNw+Om5kFdcVBVtNbSYBA19MGzVseldzzvPU+7nqf9wPNBeY7wsrKsFw3uZEXz/gln7z3m8tlztvoEP/S4YKIns4soSZJeQTRwWhtOjdD3A5fXax7Lw9lc5hJu/pJRUbKXBk8tnvcOGk5MYOk8TfAMYgk5Xe/YTQm/KN6pKttNR7ftWR4sqWyy21IoDkQxFdSrlupgRXe14LOt5xcXHd85PUHEIUy57gkg3nPaLPj4YMGfNBVPBxdDDtcDfhWoKxtTIcvNde07zy9/8RtOTo94eHbCo/fOduK+9+2FnfbGI5RDL0fd2D3aHZI/4H2g73v6vh89/VWV4B2ud6gPUGgBCZGw6uBYuoEP8Xx/2fKXj46pQg9+SNJ6Ef4oFc/WgV9cB17Soqsli4MVdV0nP6Lk4U9mmOL6D0Ngc9UzDLGPKDDksJMd4GYb/mhCCDEEEOXAwJE1VF0OhC30ntnrcoRVqQVIDFcK57vqO678gFrDomknmMSBM4TAy+2GtUZ/G18Jpqlp2gW9sdzEnszyHSiMmQ/d4GL9AzKzmdnN29ey7HOvv9Q7S/a+6nabTlsQfbedAL4WDQBQePXNFKh3PjSqzNCoEh49mD+fjiWeU5lt7Dvv3dPe6VWE/cLJrvRR3CrE5ECbRUX7zUecVd/HijJ4T1f9jvOXl6yvNzzvBpYucOo6zjYDx9ZwZC3LqqaRmICl957rMHDpB14Ez7kPXCFsbcXQNnQHB8jZMcsPHnD40WPOzs4IogyvXxPOhQ5YO8+6HxhCTWsEQkBCz0nd8KASng0DF+st5FDBOMFi3lJIsoV0N/oAKCermoeV4bjzvPQDnanpZ8Ar4ZU4fDVoCLhuYHO95ej4CJroeBddfON9CmCgamoOHpzhLy75zfU5P7vo+OtgOZAKK8lskVX63rNolI8Pl/zg5IBPn77mcmhZrzvcZqBua0xlCTakPO9azK/i+dPXfPLjX3ByfMJqdcDBqpnMy3vWfNwPSbMx86HYs/Enp89bNCuz53Y0KcX7NH0PIdB1sajRMAzpt8hgDW6I1woeiZCk/97RDoET1/OnreEHRws+PqgxwzZJ/4lRkZhHQrXiN1cdn1wNXFaHtKenLFYLrE0mld15atSqbNc9/XpAnSQGAObq+T1AipODEEMAD0U4M4YVShUUM2q0ciSBTkzAGLa5o7URA6bmfHPJVe+QumK1WMbS0WnPqwguBJ73HRsxOGMItcUuGkxtYxjgaHbYoz3NR0hivYHgB0Jw0z7ZuV33fPtX3W6A4SZcbpgG3sH2VhmAEJxYalFkj/hQ8qclwmbE27P2JVzyJR/SOzfv3cmC3+1lvG+TUe2oIrjsILSoWTw84ejPv83l+SVmeYj77Qvcs1e8vrjifL3lVef4Te9o+oFGlUYMVSIMXgMDSi/Kurb0bc1Q14SmwZwcUj96yPIb77H6xkNWD47QAPZohWkaHIZOhWvved1t6YKlrSYGYFlXHBt4GQJXg2NM3FNKxfuIULHeMZ2+0jYV7y9bztYDT9RzORYsKp7dhReACurh+mLL8MCzWCXv3nIMQnQErGuOHz3i4tlLnl9d8Mlm4LP1wLcbw9LIVBVGFILD6MA3Dmt++PiQ//r0CS9DT7fZ4q63+GWLtXUsTpMTjST1eFSlez779VPq5kccnxzz3e98xHJZpWp3e1omyElyLR3DJjgmwnQXWOZAv+umkQQFVbq+5/p6zXa7xWsk2kq0QffDwDC4mMwopavVVLFONj3HzvEBAz84XvFvT5c0YQs6MOXqT57zdcPawy8v13y66bluVxw+fo960YCJ9n9JIysdJv0QuHp1hR+ys6YdZzD/uzvXuKAVnlYDZ7XlQWNZqY/+IhoL2I5mdROJ8xjlMdr0M+eT7P+m4nzTs3WexXLF6eFBNCcI5MRIfYCng+PCWjpjCXWFtg1qDSH5PqnsH3W5coYAYSD4Pn6XuUPJbcnXbjBSO5D6o2yz46LTmZndkIVWERURfYe1AG9dA6A65Vmb0EERJyxZ5Vdw2pquFwqDW8KK7z+O8f/71yKkYkD7luoPIxzwTS2rOueMTgC8KFsDrraEh0cc1w3ywWO2z15x/dsnhKevcJcbhm2PDgPiFYvGGOfUVMDbmL6XpsYcLqlOj2k/+oDVN96jPjmCRcXGgB80MgCLBcFUDBLYYnnVeTYBjo1N2yGWBW5tRNWv/YALASsmhQO6YmOUGYJ2WkoUI8by4eGKR5dXrLoYiz9Xc9/WIsG9OL9is+k5OD6IRNYUiZFUELGIERZHh1weHHBua37WD/z356/54P0jlsbEeeWc9RrAdxw3lj9b1fzwoOE364GLoefias26qVi1J6idr5lkgGvF5nrg559+hpH/wqJp+cZHj1ks6pHlllHrEGYIWsaZQTl3IYZJ2vGuuzxoQ4KcTf0qu/l7gipOY2jfxeVVLGns3EhkfFA2fT9FA2g+bwJOofe0Q8+DYcuf18K/O2n57pGB/jJK/5nRM5oYgBW/uNjyL9dbfq2Bq8WCR2ePkXpZmAJ1tltUlb7refHiJYNPyZvG4O5ULtuEcZ1nGhZVDJ5alYUGztqaR03D0vsExwgfo8RCVJVJlTcL4iHliuSkRsJFt8W7gbO65uHqAJEuvt8YAoaN8zzpAq+p2WLQqsIsW7QSHMqQGPyMXW+yMIrVFOIbPOoGRPwogGUGKTB1kPGoyVG4s2iYP942aVMzfSpKb40TT8TfhNHW/K77Rbx1BsADqEqZluROYl5o2jIvFfgSOSpHhBKR7m4p1fyekc+XHXT3R7erbyLzkNSOnRE6azCLmsXDI44OFhy+d0K42tK/uqY7v6K7vmbYbvDe4X2I/JsQ447biuXqiOXpMc3pIeboAA5XDMuavraEKmchE6qDBXbZorVlMMJGDM8HxzqQ1K9CrvC2rGu0aXka4OUQOJWKRipQBzf2Rt5Au/MMGA18fHLE+y/XHHYdTfDEHVrYeffBS4Fg6DdbNus1fXdAa1MBmtHLOkt4QtM2NCdHbA4P+PX5S/7+2Qv+5mzF8bLGViHarb0HBPED1m95b1Hxf377m/z4p8+59I5uu2FzaZGDmsY2I0GPM1NG5zQs3dbxi1/8mv/8n/+OH/r/mY8++oDlqsHajPazRMLsbE1sz815RzewZrzrpt33Zj+7R0VV8SEkyf+a9XoTS9vm+zWGNfa9i9Uek5OuCSZmoOwG6r7jzHV8FNb87cOHfHy8wJoAfQehSBcsglYNjpofvXrGp5st63ZJdXZGfbyESgglHIDMEbjBs77ecH15hR+YSwHlROezIzIHqcRz8BxI4GFbc9bUNCEwJRxOH5WoAcCkvZsZ0BxiGKm1pq3/ertBnePIVpw0DRLWaUyGbRBedp7XA1zXFidCvWhZHR8QjOAysyM5RHcKWSt1GioKQVHMQk3vAAAgAElEQVTnx3TAavKqaowsmDbF7fjwnZVx31JLINLRWZUbsBEin9v+HoZ33/a1+ADkOiqqglETOWJy5bm5J/a+in8qU6w5RDL+pjYaFbJwoIkTllzEZX6wVWSv9J+15n80Lc0nnuVccc7EvOJiccYyVEolglQGs6qwJ0csH5xSbzvavsP1OfZaUw4TRaxAZajaJc1ygVku0KbCWUMwKWNWGkIQYlazRUNoKgZgHQy/3XZceY+aOhVsiRLmwXJJvVryvB94unGslpYm5/K/cfLKRSwIuyomeL5x0PBBDcfqqHRgInL2Zhc7NvLgHOvLNd1mS7M8nElEEHmgHFJ3eHrMcHrKi6sLPtl0/Phiw3F1yFnVIOozZxyJ2NCzbAzffXDGX531vH695mLY0G0Mm/MKWx9ixebssHF4SZWtEj3Yr697fvqTn6MqrNcbvvPtjzg5PcbYBJ8sZZbqXJlOUoyU2d3od2lG8tklwWE3hVB0Luv6nuv1mvVmE6csJhE4wQdl2w0x2i3rIlQQraDrqDrPweD5IAz8cFHzvzw45P2FRfw27r/s/IcBqXHU/Opq4J8u1vw6KOHBIcfvP8S01Z70jwJqEAXXd1xfXjFse/ApBn/ESaWupOCeVJP20mEIVGHg0AgP6pqTylAPHaMPRdJSxHOSIgCyqeUGrC1eDGvneR46AA5tRVNJTAIkCkbYDJ6Xm47rAL1YgjEsly3L40M0h3ROixuPqszj1rNvulEQHxkAUY/RVEo4p6Ge8UOR2L3jGW6/hhZpmUEn+pJhW5gfo8LvX3MUgFXBlAU3S6Ivk8hdgihxwMAYFTNZawvEc4+WcPK4OJMDYeTcZHZn8dyM8//D5AD2hu/smU9mAqgq1FqCeIbE2IoRpBLsYoGEljpolGyCH7uJJVVJS2MIJiIxLxPzNzIeCkqAyiKrFtoaJ8q1wJN+y7nzODHUktYnKIeLltViwXrT8+xqyzebQ7IdNHa4sz6jGqcUeaOa86w2vN9Yziw06jEaCPtcVGYAS6RNYX11zfXVmsOTg4Qcs2NZZgUip7k4OqA5O+H85YrfXPT846tLvrVacHRUU0sFxBKseVzWe45a4W8en/KsG3h2vuWy2/D6UuhboTWrlOCFiQkgIxxBsbx+veYnP/6UoR8Y+oHvfe87HB61VLVNzIJO602OvpeRgE/b4i7CP4ITmIKhpICVanQs23ZdJP7bbUzuI1ViQBSnyjA4+iFnZJS8EWNRpG3Pout56Aa+I8r/9uiE7x62HEgPw1CsuQGpUKnoguEfX1zwL5ueV3WNPT3i8OExWuktDEDEM/225+riMmohsupfir1T4oydfRELADlaHThuLSe1YSVKFRxSEv60L8hamRvhgSm0VQQvlhddz8swYE3NQV1jJUx5BcSyHgZebLZ0qtELoTLYVUNzuMQlor2D0cZRj/xt+mZImRZd9GcwKKPBSOZ4ZB6m/a+njTVOdpg2ybt3D4lIfrbvNJjeOgNgFBEtdsye0L59TXRHEzdDMV+25cMrO9f+lbSdzRyQiJiaCmqL76PdFgK5xPiYEVVTidAdZFiyeJFZ05S45ubrFYHKYg5WmIMFapStFZ71Ay+Gga1Cbeok5TkWleWgaTDO8+T1OcPxKtpSR++SNznzpXF7z6JWPmhr3m8sy26gwjMkZW0CSupmB9mbSCCvL6+4vLjg7PEpi6pBVGMVtiT7igaCsZhFQ3N2gn3wgGfra/7+9SV/fnLIe8uGh1UD0k3QUgXvaFzHX56teHF1wJNtz8vtls0GuvOoXWntCtPYGXKPCD0RzyCcv17z4//xMy4vLnD9wHe++xFnD09Gv4AcvXYjkuYG8Z8zRVnyy/dmD/Nd4qAEnA/0/cDF1RXrbjuq/fM93sc0wNttj45ZcNNeGQJ+7VhsOx4MG75Nzw8Pa/72mw85an1KqOSLdRYwNQM1L7eO//LsFZ862J4csDw9pD1so0o74x4t94gSnGdzdc3l+WWccznPG8CZIaS0LZQmeA78wPtty2kttCkkMAscEwMgYLO6vxiLFJ0ay4Dw2XrNCx/4oG1oqyrmOwg52sFy7XqerbuYAVCAxmBWNXbZ0tvcZxKZCt5nJmdlHJs0GqFYpzj4d5p2vTNtBqVxfyUJxAiq9TsLyK/BBGBhhJEWn7vbuH8VUJNMB583APDuVvZ1wz62kzHrj63lfaoZmVvBtDVm0eI31wh+VOdaEWwhEYzPjzgscgm7mcaKO8kPK+AVsMLicEV7uEpmAuEqCC/7WETnyEIO4RNrWdY1qyA8e/mC4YMHULdg64gUtcRuyqTOD6UeFEI0A3y4bPjWsmG13cSEQCEkIrG70pm5KIicc2yvr7m+uGCxfAgS66pr0gSMtxqhOVixevSA8+cv+OTqir97dc03lktOzxqsqWDMdx8geGTY0tYVP3h4wIvB8ezpOZuu5+l1RV+twVoWZsn/x957NkmSnPmdPxchU5Xqqmo1gxkAA7kLrOLeHo/LM57Z3Qe4L3s00mxp5O2L3QNAaGAwGIxoXSp1Zih3vxceERmZVdXdGHCxjWk+bdWVlRkZEe7h/ujn/6jAe0a8o0P6bhtQe7QU+briyaMzVosfcHl2yTe+/TVO7x3R68fooMFZ2KXu6n8ZdVWPWpmoE0ut9dn867xksV5R5CV2I+HrUkBHmZeUeYktbcsqXQ34Y/MKucoYlQXv2oK/7Ev+3YND9mOFtpnPnegq7lJBEDHOHT+/mPCr5ZrLKEUfHZIejqh7HLdy1sv3jZBfr1cs5nOKdQbEbFxZnbnYtUaagTuQ1hFbwx4l99OYAyWIbEngjA/b1IBWQjgfI9L1mnISnN42iOp22IUVfHw1Z1waTpIY5QxuucBJvxesCJgXa86ykkooH6dPQujHuEi1tyrrcQhuTpFt0BARzleauLoyQmxnSu0COTVj39rZb7OyILqs45o38o2emH9ZBeAONyDvOKi7yW0vS7dzVL0YHW2wqrFLXodNbbu6tvdvu+U6ndHaW7vx7G/0M/z9aMfp4eqmIlIIZBAQpDHFrGYqjUxs3L0dq8Kfq4Hs2VgSu870jeusc30BVjlUEhL0YgolyZRkXkmerwuuspz7QwllfbgSJEnEqJdyuZxSrNfYJERKBXZnQO1P5+k78P3iS6QpuNuPeW+QcDRd8dSWOBlSONfBiK99w905a6x8B+vlisl4wt7eABUphBI+hELd9MV6RUDHAcneiOXhEZel5efLnK9PFryX7HMY9aHMwDYY7A5siazWHMUh37sz4MIali+uIA+4nK0ohHfXqkHqQzOwEf6Aqp+TRVGVlqvLCT/577/k8nLM+19/j3ffvcfRyT5pFKJ0XUmxtShUu1Fa8b6zHbpes9aDZK3Hjyhz1lnGMs8xpcE0FSf1OayxFEVFmVdUdVObFpqgtJCX6FVOv8i4V2X8xUDx98c9vnfYI3Aloqrq3AlBWwoahBRoHi3X/OOLKz43UA2H9A/3CPpJrdlvlNcmPCsQGGOZzxbMZvOaT7nNAd1p6dKOgqscpAZOhOB+FDASjqAq0fVcNeqEVwBkXf7X8Vg1LjYESIkTkiKveD4dY40iCRNC57CzOSqR0OuxstKDbFWQyxAnJaKX4PoxRoMRts5p2uZvu8PprHass1i7Ufq3D3JbfzeOlIY1dJ0mXyJO+Ura4jytN2fj0REIhARr3+IyQG+WSLFrSd1yLB4DnnZ1bemiDTd5zelsBL+V1EktXWexZwyttuyE7/txo3Zxk3X4ZaANxLITQKAIeyml1rgWhLmTptlykg7z4vUeR/f7wid5I2KN7se4NCQvMhZC8XxdcpWVsJf6A62/v16ccDgY8GR+xXi54njQp5eqjUDYZmd03HC0T92WYDIGUcJpL+RBpPg0KyhUTIWre0Y036c78q2BFHnBYjpnMV8w0AOviDScENkmTqlAE/X7DE6PmSxzPhtf8eNZxrv9gr8b7PtmMWUFpnHFGAQ5kYJ3ewH/9rDHar3AzAtE5rjA+na5QhOkIUILb323DMeXK3qoYQ+vO5+u+eR3T5hOlzx78oL33n+HBw9O2R+NSNMIqVW9tG2n/N8Lwub1VvyzBfdxNYCMpSor8iIjLwrysvSldK0iIdqcAFNYyqykLM1GBhrj0f8Kg84K+sWa02rJn4eSv98f8Jf7fYbC+Li/6YoZ5fNNgojPloYfTJb8JKuYRn3iowOSvT4qUNuGhtvUsjkc6/Wa6XTOepHtWPhdBRJuXOG1nqCtow+8G8XcVYKhswTOhxeF8AnPggqEt9699LTbCqarQw9SUVnLOsu4ypYEUtMPIyIELi/BWFw64qqUPCktZ86yUgIjIein6F5KpTzU98tFzq63x5dlW1fhnAGnb3Br3zwTbcv2G5T/LyNteTpuTOLs8Bxh/ycSIHi96HWsdk/bGntDkiYEcH0+X3buTa/mpqFto3Ff/1b38X1ZaXfUzUw4IRCBJuqlrMMQVF7HHLnFZbw5w2beXqIoNY/UAdK7gnWkUf0YBjHFfMFcaM4LyzgzOKfbGnZhoacDjvt9pHNcLhYsqkNSFXU25A3PdOtPn9MgnEDLkMNU87V+zC+XCxbSsu4It01ddvNb1EzaK6e2smTLNePxmCiNiVQXhnbjdkVKdBzSOzxgdrVgssr4Vbbm4WTNu0cHnMiQUBYIW2e0Y8GVCAMDLfigH1Lc2WdaTiErcSvLBEGhNII+QRIhQnFtrP6OvfLigPWy4Gl2zng8Y3w548WLSx4+uM/p8SF7o75vk6sF1npBsJmKWkluAYSctxKtw1hDZUrfPjevKMqc0lSYjoLghb8/b1k4qqygKqu6ctMrPa4ykJeovCTNCo6rjO/Ikr8/OuQvjnqcxtqX/FXdUI/ASQkqZGklv5zM+Ofpis9liNkfMToaEaSRf2Q7IajGyLfWsZgtWc1WVHldCupuE2FdX+JmcSnn0f+GQvCVXsIdHD1nUV0QKvDJe5I6b6UZx7ZVDR79Ly8d49WKlcnpJz36QYQWCmcLbGZwRnJeWR4VljHec2a1JBn00L2kbQu86we7eUzd8VhcxzMhbjjidqqt3l1v75edmdbkts2kmmxr9Dj3llYB3AEKJ1/RAvDV5L0ACg84cvMmvUmwXTvAiZrB3S6o3oZYVjtXHdlhhUChCXo9wl5CtVrhqvJmBnCbnBXi5Y+59t60JUlaEaQJatCn0mPmMuBFWXK+LskLR9zJlu9pxXGaMAAulgvmZckdqWo3trj1efr76jLcCkHFYRzynf0ePzgbc+kM012m3DA1L8mbWWoPKbKc8xeXDPf20WGAkg1EcZMM6L8qpSJMUwYnd1gsV3x+VvDP0xWnz8f878d9jlSIciW4OrPdWV9ejmCoE/7yzh7rShCcjRHLnI9XlnMcubGwPyLAQ7/Wzod2/TadA/3b0ru75xnz+ac8fvKMz04f8879ezx4cJfjOweMRn2U1pSFbXCTaHEC6/hwVVVY46hK37SnKAuKMsdWtWIkm1JA/03rBNY4ytJQZBVVXuJqjVwaB6XB5CV6vaaXF5yWBd8WJf/XQZ//4/4BdxMJVQ5FtfVYPFZ+gAtiPr1a8MOzCb9cl4z7Q/buHxPuD3yyJBvcD4FHNnBO4KylzC2T8Yz1MvceGAK2yv9uXOBsPJPOEVpLHzjUkncGKfvC5wOoxtSQBmFqxVOwif/TXWuN4qhARszKjGezFdYZDtIefR2ihcNJReUgK+HxOuNxVjGVIbnWuDgk7PdRSbpRAF7qk9/ewH5Idct1Nmu40SC6Yezd/S3YOGW//JzzNtoRcJ1wgOAtRwKs6feegK79tQ1vLrYyzrvUukJf393w1pIvBevgyzuBkxCFIfFwwGqxoMqyJvndz3+zsLuPs7E26rfU68y9ED4soxQqSUmGI+bqBatAcJYbnmQlZ+uSd3ohKM9AA2nZCyWnKmRuCmZlQWUhlE0tutw6vyfDtpvOeYjhqmRfB3wwiHkvlHxa5WgX1la+ZCMIxLYZ1TaOEdjSsJ4umVxOiZOYNNCtddlcyvMAhwokB8f7sJyzXmd8OJ7yD4+e8jC8R7ofMggicMa7uJ2qZUQFLidSkv/tdJ/YWrS9wmY5Zi0Yl4K1kVRFj3gQo6O6cRAb1/3OpHvsDSHJM8vvfveYJ58/Z3844Pj4kHce3mV0sM94PGe9rigri3Te2q+cpTKGIvcWfFlWlMZgaBLMamWp2bVS4KykKh1VaSiKylv+TiJtXXJWGtw6R2cZe3nOqcn4trL8+72U//trDxgEBlWtqTvzdCYVEBKrAqal4r8+uuBHs4yrdIg6PqB39w4yCXAS5BbCXm1IOIcpDfPJktnVgjKzbIS/3Ixhl4l0OZgD5SyJtRwIuJeEHCchqVkTOI8LsOkr7t3/KFWXADawPM356/CEUFgZMC6WPJ4tiJ3iTpIy0BrpSoxUlErzJCv43WTFk6xgJgPWQmDTGNVLkFFAJajBfF7XeveDcw0CUY0r0XrznPO4AtzMV1tu0AkBXEv7+rLTTfPSyn9wzu0wzTeH/gg4ADc0KbuBtpTsmplsdPeuI++LSvcdp5a4+Uy3nf2NfHr/I6idDv/P6oBwMKTozyhXK2xhfXaw6ygBX2AytjLkoc3NCOKY/v4e8ziiLBzLQvO8MHw+X/HO6ACc8S5yZ0mU5CuHR/xoesmzdca9Vc5ppLme43xTDLfJvnZgPQzwfqj4zl6fn1xWPLUlmQqoml4DTUB8S/bUykGj6BvL+GJMf9AniiJU1DTubVaaH7OQAhVKBncOqFYZ4yznw+WU//LkOX11h2+OEsKgjgubWotwDuEMwuZEGv7sZIiIFcGLCdF0zael5HwKeVmwLhLCvR5REiGl2HaS7TyrxiaWaIyByXTBYrnm6ZPn6DAAITGVozIeFc5Yi7EWi8VZV6Pvui01w4jawhbehrRWUBWOLCuoigpjDMI6ROXAOkRRobKcYLViWBY8sAXfCgV/f7DHf3jniEFoUVWGqEq2YuVSglYYpZkY+E+fPeGflhlPghAODzl4+NAn/gUKxCalc2M8+NPl65KLZ+cUrfXfrKHaMr8JEKkxc2sNTztHYkuOAninHzFUjqCyHiIbao5VASVo4e9J4hW9VunuXEJKVsZxnmWcFQUj2edAJaRCIh1UQrDSIc+Lis9XOS9Kw0oHGCUIDvZQ/RSh5XVYFfea29U5/3yt62yn3X10fV7ErZ/Bl5hrvpy2pszJtxoIqC0C3A6L3UjNIb4kr62e3WoQ1hy3S6Lzwc0XaDZ3Y/1uH+XqXgA3PSrxupvoT4SaufIYOqI17H0PFIHqJwSjIflihamWSGPrDqY3o1pIdgztW6nDXIVHGyPW6FGKGMbYdUEm4Vme87vpnL97eIwUGuEqMCWR0Dw82OOniznPZkue9ZecHve9YGjc5zSCu7nTRlpv3EPCgTSWvlR892DE/eklj8uCtQ1YSp8rsu1D7b5WG77oYD1fMbuakaQpA91Dqu0WO64Zs3SEg4T0ZJ9qveZZvuKfFjn7FwsCpfnaMCYIHLh8U+fuAFshjGMYhHx7LyUUij055R9nOb8uVrywJUtbsLQFpt8jTCJUECCUREgP6dLeekcHltILvNI6yty3IUasEUIia7AaVcfvbX0WIUC5pnvAZl5cjRznHBjjKAtDkVeUhW8x66xDGIstC2RRoYqKNCs4yNe8j+H7Pc2/2R/wl3cG3ItBlStElW8ycoV/bgQSowIuK8FPxwv+4WLGh06xPtgnuXuH9GCIClQ94iZsI9ol4SzkWcn0asb0cuq9EltNf25KVG7WT+Pe8b+VtfRdxUmgud8LSV1VW/+uPV5gvcAPFIQdBbQ5X/daQcjFuuTxMmMqHO+kQ4ZKEdUJhRWauQh4luU8LwxTp8hUgNOS5GAPnSY4eS3jYcO7toa1LdS9Z4TNvbUm28byF+0cNVe4Hoq1re3/xhq8vzddL2tmJxGw+2L7WOdjzsJa+7KGGv+q9EdoBiQb0fJ6x+O3oaTBV2tggK2PUu249ej81VUC/Bu+a1tT694whI0CsK2/3uio+aIOhzeUunPVjfg1/6wAFQUEwwHhYs1qVSBticea656jYWTQVQxeN4dCAE4ITCBx/Rh5tIeZrMgVnJWGj1crxhUMhSQUeKtdCg5GKWmU8mKVcb6Y444HCKU30MRb90XndS28cV7LM4ZEad7b6/O1dM4ns4q5ySmkppA3VE1vAcQ0qG2+i9x0PCPupcRJSJQENAmHDurEcx8DlqEk3R9gsiNm6xWfjCf842RFqhSp3uNhv+97YFXlNkaAMQgMezLiO3spfaWJghnJbMWHZc6jdcmkysnzHNvrEyQJOopRoURoUVea7TCnjpLkmgQCwGF9X3gBts6abyrkdldP854DKuMb+1RFRZFXmML6JFJjEaaCokTkK6KiYFAZTozhfWn4u2HC3x70+cZ+ykmioFj6uL+raDvjCUApbBByWQp+Pl3zn59f8ZPScjk6ILp7Qnp8QJAErQK/lZpae7BsCcv5ivH5Ffk6A9tx+XdUto2+13X/NAqAF+qhLTmU8CAKuBsGxNUS1eq3/njhrFcClK5xondNmeYWJQQhZxdzns3XVCLkcDigLyF0HsuikIqFini6XnBZWVZSUQUa4oBkb4hOohqQavvU3Z/tBdD5JTxE+gYDYMc5ceOXbhrHl5MaJaCthrnGXG4Q/nUyrXFW1grAG0n/ogqAMUYgN+GQ16Xt7djs6KYn+u8hk52HtWw2pWhFXvdKby95Ibz9nsUilUD3UuK9EcV8TTWdeUbunI+rOvfagv4atVNe441rgeuFRCeHZE8uKJRkIiWPreWzdcHXE0mIQrgKgSOIY/bTAc9WK2b5krI0hDpsKxa8l6Fjwd+oe3rmrHHsxRHf3BvwYTbhMitZWkvRNkO5ccbYhBT8n8vFisnllH6vRxiFdafCRmh0vy7QcUTv6BBTVsyN41eTKcnVglRr4uSEw7CHFmuoSm891oiM1I2XEiX52l6KDgOGoeLOdMGP1zmfrkuuytIL36RCp5YwjdGRrq1PiZD22j25VgVsdkZjwzoM3eCb1+Pb42qN2Tnh8wNKS1EaqtLgSgOV8spMaXBlgSxWJPmK/argAY5vBJq/6vf4u7v7fL2f0FcVVCuPjbAVRRYe7CeMWRDyi9mC//Jiyj9O1jxPB0Snp6Snx0SDFKd2PFGuI7As5Ouc+dWc2dWsvkRX+Btusmo3Jgk08XvlLLEtuRsr3otD7gCxrfNfWsbluwSi8Ml/srt2OmMTHvwHqbhar5hkOYGM2U9TesIR1J0jCyGYS83TrGJiHEUgcKGCvQHBIEVE+tpSv32HbvM9nyDp70VcO+5LLNlfg66BIHVTjWhWj63DX9uqgbVOGJxw7i1VAODWvNrbSQh3zT1Wu6Ouu7JuOUXzU2vkyvl63aYN9wa+5iUtZHfO9+Wlri9E0KhrsrYsXFYyznLKqgDj0M6ihGmOrmnXZrjxMuzaIlZCiUOlAb2TA4pBQnEVMMtDnhvHrycLHgR9hqLpoOaQUnBvf8Cj5ZjFOuNiuuDe6X4NEdtY6Q3T7jb42XFd1rkACvizw31+O1vxPMsYW8MC4/0d7a2KnXM0Q67Bf0rDYjrn8uKK/iAlSOpmRk0pkFMbF6twhL2I4d1j1kXFhRX8cDajPJtjgoT/cNJnXwsC1mCyjtHowJVgBBrH+2nI3ftHfG0Q8+Dsih9MVnxUWZ4vC2bZknxeksch8bCHTkNEonAanGosGdH2FfDmfjOuBg63FojNc2vq+lvUP4epLKVxFEXhE/0qBxZkJRGFhapCFhlBuaJfrblrSt6Rhu8nIf/2aMRfnxwxjCTalN7qNwXtjTTJmEpjdUQuevxssuI/Ppvzj+OST5MD5MkRw4d3SfYGoBXXAlT1nAsrMIVlejllfD7GFNW261Y0IZddPt0R/rXWI60lMQX7GN5JY95NIvYqQ2RAO+nj/024wBqIQ+8BaE4Hm3UpfOkfQUSRlVyt56xMxX4yYk8LUlMhbUUlJQshODPwwjhmCColEZFG3z1CDhKclvVq8xd5nWTcrn+jfe7Nzyu43s0Jf2+snPsfSG08pO3a2GAh2K1pE60D6e1OApQSxOsnQQjwMUO6+ueO1vya5LWzjsXTxvB+j9O8hmz7k6KXjKVxE1sESIlMIqKjfdKiIj8bY1cZxlZ1PsAN7sybLnDL9Zq3jQCnBeEwQe4NKc8mrLKSs8rwi4s5f9uPuJNKpJTgKgSW+4OEkzjk7PKK31xccnx6hNIBwpraE9D1BrAVz9y6AeOQpuBBmvCdfsqny5JHecbUBhQCbFcJ2IIbbl446mJzirxicjkhiWNO7t0hSHxLY+dsZw033dwkKo0Y3T9h4uDSOX46W2AfP0dXI/7qcMj9JCJsFA5bbISZK/CCqCLRAR/sxYx6p7w3WfOj8ZpfLwoeFxkXZckszyjWGUUSYGOFizUiClBhiNKqzhOoO745nzPQxMFatbC+5VboG4M1TYy/pDTG4/tXFiqLMA5VQFwZYmPomYw9m3FKxTcizZ8fHfD9gz7vpQF9bVFlgTCF9887S1vPiAatMTpg4UJ+djnn/3l8wT8tS57EPdzxMYfvPyDaG6CCusmQcBulDFeHsj1s8uxqwuWLC5bTBvWvKR9tyvI6qIi7lSP1OhLWElUVo6rgYah4Lwk5DQS9Mke7OkTmRN3REP+8ta7x/3fd5/X8SgVBwidPr3g+n6FCxZ3BgCGC2PqkwkxIFig+X645t465lJRKopKI3ukhpGELdrYBhap/v9JT10nnbP20u2GA12GYb6R8+4Npd/68suS6f3Xe73wPPP6dEMLpt7gMsMuCX0Wi+9s1AbVdCfzqxdh64kS9rbe8/p2M9rea/Lz6uN/OQkZ6l5YWyH5K//QIgSO/HGNWFlF6y1m6jaK2WwZoO+6w29Dnm6s5KZFJSGeLHfEAACAASURBVHQwwvQS8umaMY5P5kueLgacRAkDrX1CnCsYhTEPkpRLOeXD9ZJvFoZDqXwHQbocsIMI2MLe1tLMWaBEVGvSUPPBXsyn64Kfn68YG4NTggLXQiJvmUtbSkCd820s62XG2YtznxAoB+hI+cvIOqul8Z0rkEqTjno4e8zcOi6N4+eLGeGLMSsH/8vhgPeSCB0AhUPQhAMc2AIhDMpYejrgYaIZBinvphEfTzN+O8/4aFnwaVFwluVMS80y02ShItcBMlSoIEAG2renVRIpa2jlbiKZA9+r122Ef1lhqhJTlJjS5+UI4THxpbFExjKoHHum4hDDfWV4L9V8o5/ynX7K8TDlKNb0qLzFX1Zsl2vWXR5VRKVDxhZ+Np7zH59e8v8tSh5HKe7ogMN37tHbG6CCoLXOBR5i2uHBo5ooTLbOOD+/ZD6dYsuqtnZ38rIap2ATQmomoOk26UA6S2pKTm3BN/sj3o0CRq4iMiXa0iIlNjkHqBB0WF+rUTS6yqnEyQAjY359dcF0nbHX2+MkjUmtJXAgUFQiYOYkH40nvLCWpRKUkSIYJsQHQ2yoMBIqWefwdMa1G7/e3n1dQSY82JqTbTvgdvytcrRJrHzrSv0aaqfR56NZ6XBOXhNyHgRLgnXCFW+pAmCMEVrT2VC307bw76iy+JabonnNK4T39lOgqSRwnY8F3K4EtEhm3dO9sc/vD6BubKv7/gYeGQkuUAR7fVLfK5VcOKqFh2/1eOeuhQJt5morc1bUF7iRAXWEtdIk+3sU/R6lnjItLM9Ly+9ma94bRPTDAIFHzQul5f6gx6eDHr9YLflkPGOwnxIItblOd0zipjecF6i2RJo193oBH4wS3p2sOS9zKiEwUlI5aJvBbMyqzoDrFeXw9eXTOWcvLhCBpq/6SF3DGXddq8LPmwoUvVEfYWBq4OKJ4YerOcXFDGsM8qjHO70QHQgwBYLaSq5hgzEO4UpCJ7mjIo4GAffiHh8MIz5bFHy4yPjNMudxWfGiqBgXgrkQGCUwyrd+NlphlQQZIZSuMeSpBZ7DGYszXgFw1nhEPmsIKkNsLU2tjsYRO8vQWU4E3A8l78aab/VSvt6PuNuPuBsoFM4Lflt6F3mTuyEEoHBCgQqwQcJ55fjFdMF/fnrOf5tmPE8HiOMjRndP2Luzjww6ShVtf8LWdnDWURQVZ2eXTK6m5FlFq7Q1pZ7tWmjOc4PCV1vzoTWMqHgvEHy7H3MvEKSm8H0Kulpwo3hGsfcAyOa9xvtYrycpqYTmInP8drXCILkfpdwJAuKyQFqBVYo1ksvS8OlyzpVUZEpBEqL2h4T9HmUgKSVU9fLyYdebGnPt7onNEAXUOBJiwxu7zpDuWv8yssPXpcaRI7xyZdnE/l37H2wwJSRvMRDQId6Eus1dfAM1zcrbv30dgEc1a8T5q+fT0ZEFYvPj0cBuFkjd64rme79nxOCNp5sG4m56WVdPCLBKEu6P/N5XkGMxqxWuNEjn2k6K0m3OsFHaatWtkzjovTN+chsL2whBMOqjRwOyOGKdGSYEfDRf8+dZn7uDBO2UF4SqYr+fcDTok09mfPTigg/69+kpDUKzsSh3tMHuBLQM3iFMQT8IeHcQ8+fDmEfnczKryIWiql382xxTbHelatxNDmxpuTi/IogTVBiQ9iNQm1JLf3i9joVDhZLewQAhBFe25PK54GerOZxPsFXJvzs54LQfkQQaLTMocy/8gQ14kANrECLkIIo4SBLeHfV4b1XywWTJo2XG51nJ06LkrCxZZJa5M6yQrKUkk4pCRFQywEqxkYnOPzcfknO+Wt5CiCVxlsRWhM4Q4aGLD5TgWHvB/04/5Z1BzPuDmJNYg7CQ5zWmfwOE02wun6SIFLggwKqYi0ry3y+n/LfzK/7fyYInaR+O77D/8B6jowOCRFO1SliD7rk5LU5Q5RWLyZznT8894p/FL2ChNkrpS2Rk+5l1KGd83b+wfGuY8G6s2MMQmBKo6meq2qUltYA0rrP/O+h/TWJSjf2fOcWvr2Y8qUr2ooTjKOFASELnEEgKoZlYeJHnXFQ5i8jj/etBTHS0h4wDrMJ77L5wYm7jp60rQZxrG0W9bHreRmq3vPPgScqZzSNt+cDGnBVCeJypN5TeMCTAxpq6rjA0EL7tRn8NcoCTm2ZABod9xSZp+9z8Hnf9p0Uv29INdBVbbgEnwGpJuD9ER5ooCVicXVDNlr5JSWXQrXytBXv3cjfMo2Gj6wkpkM63B5aH+4jRGLMomAURH6/XfLYq+EqVcCAVlA5cSRjEjJKEAZJPL1+wOjlib9hD6QhMSVNMumXGXLuPminbCukq7vVi/tfTER9dXbCwBSuhqYSovQCdGDHN/HQ0RASgwRmqrOLi7AIRSk6jI0JV16Y33hIsCN/WVgiBDCX9wz5R/C4vAsnkheTHsxnTiyVPMsP/+eCQ94chezomcPhM+a515+o943IoSpAZidB8tRfxXn9IVQ3rGvM1j6YLXqxWPMlzzi2MnWbiHDMDa2Ux1is8QtSWoHWt0qyAwDp6wrInKg51xb60HKuAk17M/V7Eg37Mg15KGnrmqMh9aZ81NehOI6g3uPPoAI+Ep8hlyGUO//DsnP96MeGXRcXT3gH69JCD994lPRihggBzEyyd862rnQVTGBaTJc8enbEar2uWcjuU+O37QiJcRWwsI2O4F8CfHe5xSklqSg/j3Coixsf/pYQwgEiDqNg0/2lQAAVIjRWKZWH4yeMnjPOSBwcHHCURA1cQgE/+0wEvsoLPl2vWBBRIbKBIRj0GR77dcTOTr8OurnkFROPckkipaEoB/UeSDpLE/yQANv1oGqNHOYFyog51emXWuVqpfcMTI/9YCsCr6Yb9J/CMSCJooixCiNt6+dxKzXkE0msEt3gkrp32S6v+doMiO4KtS0LU2O1ukxPQS0m0Jur1yK+mZOMJ5WJJkZeoGgFVWNf4w7av2LGkLd7qd8JbG0JpQh0TvXNKcTmlPDtnVgkeG8GvFhnvL2MO9oLafW6Q1nIn7fG107v8+MknPLqa0Isj9nshwmqg2haS7aV33R11tntV0Qst7w9j/na/z/NpzsQpMgfG6TrBjE1I49qUNYqBVwLyxYLxC1DacXJ6RBhqv/TEBqtdddzXBALdTzj8ykOWacrq2Rm/GU9YLlYsf7fmb49H/PnhkHtRShgqpKkREq2pPQE+pwEhwFQIodBVCVIRCM1prNiPUj7YS8mriqui5LISnJeO87LiMrdMK0tWGayz9V5xNUPz9xlqSaQ0B6HmJFQcB4qjUHAUBiRaEkpDLA0hObIyiCaxjzpVujmX35DeEpcKpyMqoZmVjk8nS/7h8Rk/zEs+FgGT0QHR3WOGD06IRgNEGLTQtJsHUuNYOr/Hy8qyGC84f3rB9HyKMx3wpps8Qe2SqJsCtYc5cJbQWfat4b1A891hn4dBwKgsiIzZAP/USo0ElJbQeD1ofhybigIBQURuJefzGZ8uXhC7iCOdsickYVV58B8dMBWaJ2XGo3XOWgZYrWHYRx+M0IOUsvHY1LfbLslaiXsV+btXCKl9Dkgbqtp86qei9uzdyny/lNbSzbS1/evqk92cks2xDRN9I+nNUQDgOsNuqNFInW9K8sXkcut/vZFkm7m7zSsaXvXlou0BXct07bhHXYejOCxO+6YlYaDRYUTQSynmc/LlGrPKsXmJKyuEqbuLuToeKsAJ0RTG4aTAagGBRocBOkyIoz694R5yvuTsk09ZlBkvSsmHq4w/W6z47miIUtrXxGM4jCO+dbDP46ef8Wg84WhvxLA3RCtZu8Z3ht2GKBqBtPF2CEp0lXOoAv7tyT6/zi+5WBcsraAUHont+rlumM6aP9rKsJrNudKgleTgYESYBHVmeh27dpvSVoFAaEU8SvFhcMU60jw6P6fMVlydz3mWGb63N+Drw5ihkoSiQIoSXEHbTAjYhECcBxGSllBKQqHoa49Kd5hEPHSCzAhW1pFZR2EsVeWR+6CTu1Dfo9QCLRWRkqRKkgqIhSNRohaExt+LrWpgpl1kvdr6rd3wTgYYFVJYxZOs5OeTJT+6mvPP84KncURxsE94fETv7h3ivQEi0G0Yr1UnOuEXV7uUFuMl58/HTC5mVJnzShl4r4tovt2EAdiEAmrQpk0Y0iJsRc+WnLiSb0QR3x32OLSW1FgCC5v0L1fjZIBQAkKN7+dg/LhFs+YAEWBlzHhd8fH5FZnJuT+8w3EU03OO0PiAQik15wY+LwxPKsNShxgt0QdD1NE+LokwNb5AB/fwC5BASIVUHsi4bQ/eKi3NGLv05UP9u4lEGybyY5QdttJ4ABrX/1btRL2n33oPgFSusdlvIbc1oS876iY96vWVgVcv1Obxic7fr7qvPzlyN4xqZ4BNJ7ktcwKvzFqkz6EKBKLvgW/UoIfOcqplhl2ssVmBLcq6e1zT6tafT0iBkwIdBIgoRCURYZIQxwlRlJIclNirMeNfHJJPZ4xLzadFzu9mKy4OfPkfrkBgSRXcTyK+ng55vF7zeL7gYJhwFNVx3m6M9ybLxXV+2wrKjDiwvHfQ43uzjCfVkkmRkwvFQgY7YC7dbiu1FdZqkJ5LmKJiMZ7iURQdo0OvBEjpBZBsb6v+ngSEJBwkKK3QUcAyDnl+dsliueTF1ZInq5K/XvX4xrDP/VjT0xKJRDoJVnXczZ2xGeMFsqhr/6UkloJY+AoAlKjHJryHrMH9bZSkZus0w3e118HVaH9NK2MM3vNSf94mQokarhmP6CdCnNAUVnOZ+b4PP50t+cF8zYe54/lghLhzRHJySO9oQDToIYINyt8mft/Mt89XMZUjX6w5f3bB5GxCvqrYxvnvNuHpzM8ua+gI/8hUDKuSr0SCb/dC3g81vXJFZB3aNS5fQBg/WiU88JJyXgFoPABtGEmAillZxbPlgo+nE2KneDgYcRQERKZCOkclBUspeLoqeZSXXAhFFmhcrIkO99AHIyqtsHXGXgPQvLu0t9/dKHSua0gJ4cNwSm3tiQZ47aUccJcB/ykwyz/gnreWitts+VvOX6tR+o2dlT8KEJB8xfC3FuJtx9QWpBNii29vfb9Du+fxSRqvxiPsJtK82brbvyzd6BWg7s0gJA6DUAohJSIMCAd94j2DWxXYrKAqCopaCcBanPV1WUIBShJEISpKCOIYHcXe+hASwor0wQnD9x9y8bvPWVaOszV8tMr4aLLk5MGBF2bWl5GlKuCbx8d88uRzPplOOehHHJ30QUUbYdgqM7dpkF5BEa5EGEGcxHzvYMCnyzUv8oJlpVmpwCs/AnA7AFKtTtUIpY2FafKK6cUEJSRCKEaHQ4IoQEkQom4T20Ly1qeRCp0m9IOQIE1YRgnz80s+Gk+4mC/5ZLbg3xzm/MV+n4f9mMMkZqRDL3BMUc9PkyjYnNR5odx4pJv5cPX1tzibqI/X9ZudJLYmstOctwXPsdQ4xlxH8tMeDEcqkAEZAZPCcbYo+OV0wQ+uJvw6L3miQ9ajfdTJEYN7J6R7PXSkOpED0VmbTXhCYJ2vwMiWOWdPLrl4fkGxKrxC5H3hnQd1myHQjMfPlW/3axhUBacYPuilfL0XceRKIluha1vZ5wj48WsBItQe+78V/p1wo5MgNMiI83XF7+ZLnpcFR0GPe3HESIK2FiMcuZJcWcdn6zWPi4q5jsi1QuwNie8coId9KrkLxNM88s34XsXvRK3gSemxNmqHWLs0WuTHL58b9Pekm03NrXe7e6rmKw63yYd+A+mNSAJsvXjuhoi06PoIrtNtzXtuuoHtKM3NMZtO9eGXnL7IQDfzZVFIIesODYAUKKWRQYjsOwLn0M5hrbcSXZ301VigUnmB6IT2HfgAhSEMBNHhiKP3H3DRiyhKmBWKz7OcX4/n/PW9O4RCISnB5MRS8PDOPoPzCy4XK56OZ3z7YEAYxLVrvFM/v2XudQN5buMhcAZpC77eD/n+IOXRynBRFEysJhch9qY+Abu+V+G7Ajboha60XJ1NEWiEk4wORwSxqmPZrhNyrZ2ItTwmUMSDHkkQseylzJKEZ+eXXC3mPJ8u+eVqzXeHMX95OOQ7gx5REBBqhRIVwpTeOheCFmCnazVv3X9jodrO1DTzJdnEspuBNv5y1XmvqXVvLH5Re2E0ToQ4pSlkRGEkj9aGn01W/PD8ig/XJU+VYN4b4fZGpKfHDI8P0WmM0GprXr2TpeMvdL7tsC0Ny/mKq/Mxz5+dUa6LVpBvh3s6OQgtye0t4LzCo5yhZwx3TMEH/Zhv9hLua0irNcp57IJuMpi2zrv9w8Bz1SY5kHpOG3wDEWCd4vOrMR+PF1Qy4sHwgCMpSJ1BYqmEYK01T7OcR9mKc2NYRhGlhuTkDuH+EBkqqlvCzm0/BHfjx1vz6Z+0ACVRStVrsYFcf9m3Nz6H5qg/lWTBLWfWH3qi9gQvOdvbngPwKkt6ax5ramp6Peu5/TE1JbW3kmMrH03sfviSm7o1efxLQTfN+kuOFt26Yi9MPH64jxs2MUPTuIzZyJsWGrXxmQlR1yxLnNuARTsnKaREhAo76MH+CLcas5aaZ2XBL1YFv5gu+aAnGUjpk+CEIYhDvnJ0zOL8Oc+Xcz6/mvP+vSOEcB7dsEGE2RX8N7rvLFQFsRR8az/hSWE4v1qzKHKuAslKC1+r3v3ylnXUvN70CgCHqxyTy7mv2HOG/eMRKhBItW2Rbrxa9b1riUgikjtHyDRluTdidXHBo8mUabbiyWTBbxdLvpXGfDDs8X4/YS8KiXSEdhZtfUMaQeWt0gZDgI6U2Koo6DKybu16c3f1H6JxqQNoWnAdUTsOUBghqAgoKlitDZ+u5nwyW/GrZcFHueUTA9O0T3UwItzfIz0YEY96BHHQnqs7J9toegJhFVVhmM8WXDw/5/z5BeW66kBC71IjMe1NDKf27Biks8S24oCSrwaS7+71eTfSDE1JaDzqn6jnTjiHxPrpiMK6FXGnh0NzbiFq2N8+i5XhyWzBxbqgFwx4uLfPnoDIVgjhKKTmSio+XS94WlRMhGStgEjROzkg6KcYVcfpdy3z17T+RceTCnhPnpK1MijrRFVRb/XdM91gOL3kWn/y1BnurjHqFGCbzo9bkqjdVU0Gyr/kLX5R+iMoAAr7ChyAazOzZQZ1DmgEyY5VsLv6uixVOA/EJlwDKNRE7bbNtqYdcPd6XeXujXx6fxB90S3bnZxaigpRW2Y1U6mD242nWNj689okcdfO58/jEBghKLSm6qUED+9RTXKKRc5lGfDbouRHZxNO7u/TCwPfmMhapDJ87XCPyXLOs8klv7m84uTOHVIR1H0LGobvthfMNeaJZ+qmQinJvUjxvVHCeWGZXmUYU1AJRa6axMbbVkV3ITVZ5ZIqr5iOZzhXYWzJ8GBAkkQeLEiI7UUmvAXme2kKpAyIdR8ZB0TDhPXlgOVkzKfzORerJR/PVryzLHkvybjfSzhNYk6TgNMwJFEOLRQK6feANRudyDWue3ODJl0/m/btDiZCK3y8Ze1EiBMKKwRGCionuSwrXmQlz5YZTxYrfrsqeFxYXqCZhAmr/T7B0T7Dw33CuoeCaqoltpTv2pJurH4HwjpMaZheTrk4v2R8MaZY57SlFtSLry3Fcp057poktZZa+76Vs0S2ZGQKHkjL94c9vtXTHCtHXJUo6lh/s56cR2kUWkEUeKCErvBv503iVICRCR+PX/BkucJKyclgxFEYkJoC7SyVkKyl5qkR/HZV8txallphY4U4PSA8GiLS6KU1//I1DZcGU8X3I1IorW/uiPoS+oOt6H8F+kPuuW3v3VK9pq5Z+a4O8VnBWw0FfK0Rgv9TdObEywWx+RixxYs2rqpt2tUPbqKGBTTusOu21uavBizI30KDiOZuDCn86dPG1qT1orzCetit8cc/ty44UzdpdgtGtyM4uvocO2ezQmJ1gBj26T98wOLphGK2YloUPCorfnQ15bvDmL2DlH4QQVkirOE4TXlv2Ge+mPHZfM7Dyxlf3e+RqLpHgGsUgY3ScuMgnQMqRAU9GfNeGvA3o4TLvGKdGXJTYVBUQraKznVQmc5KE01TIm95VnnBdFxQmYKiKDg82iftp4hA0lQYd/M0W5+LdIhQEgUxYRISpjHZ3oBivmAynTCezPlssebns5yTZcXdaMW7keJrScSdSHKYKEaRpicFkQzr9q+A810ekSXCemWgtQ0bYbqjtLlGkRN1vbMLMVaTGcGsNFzlGRdFxed5xmdZyaOs4HFRcO4EWTKA0T56b5/e3pB41CfqRRAInHTtPkQ0GfYb4QzeC2UNVHnJ7GrJ+fNzJlcziizfTFzrFmx3/+b9NrmxmeB6gdbzEFrLsCq5Jy3f6kV8f7/HQ+UY2oLAGpRrBKythb9FSAdJCEFzv9eFPzKgFCFXueWnkzGXWcEw7XNv0KfvDIGrAMilYiwUHy9zPi0sVwiKQCL6Mb33H6BGPWwgt0Kf7UtxC0zatXLYLhe0CKlRWiK0bPsJdBWMXeyALY/AGyvaXkJ/0D1va1e3iYbG+yiFu0EGvjn0L64AWNU1LLqa+QZycmsSb1qrtbly7dhXUa2seaS6jd53k/fv7U5yaealFuIvO7Kz8Bur/7ZT7gKt7fak3yYvaKyQEAQEgz7pyQHF6RHrywmL9ZoXVvKb1YpfjOfc6yf0e7Evc7MVYWB4MBpwthzx4/MzfvbsGffSrxBHPlHRO6FuZ4T+nt3GGqREKMVBqPnOIGBWpVydr1iWJaUVLKTwzYIa9+7WQLvzsvFwNNcwhWF2OaPIS1xlOTwWpMMUHYqNk0IILK5OyN9sFOEEQiiiYY+gn1Id7JEt9lmOZyyvpiznS16s13y0zhjOVtxVgnta8c4g4W4v5TgM2Ati4igkVIIQL7cCERAoh5agmv3mQDiJrcM9xvl+AJWxlDhK58itI6scqzxjnFU8W+V8vljyWbbmua0YS80qDFn1+5jBkHjviOTggGQ4Ikxjny0v/Eh3l1OLmNh5dLa05OuSyXjOi0dnLKZzTGU689wcfJM344Y1UD8TgUNbS880JX+K749S3o8kB8WatCoIXFX3v6j3ibNI6ZCBgiSGtl/DzhqTGmRIZhU/v5jyq8UUJxV3kwF3k5CwWICzFEIyFYpnxvGr2YJnxjHXijIJUXt9Rg/vQi+pk/86Y9xN2L1h1DdRyxG1RAQKp2QNllYrec0ZvpQe0C9Iv+dE3Fy79ubQvwIOgHfJNdv1lTH8dpnajtvxdUi0V9s619bi7nwibmQN7ffafIAvlaKw6QbfdbbePkI/CRY6lvz1WROdw3cfWYMrtuvx8Z4FgZPgIo3rRZSxJjk9wjy/IJ/NmZuSF2XIT8YrvrlXcJrEREKCyREmYy8JuDca8dHVlEeTM8bTA3r7A2KtwdVJca01/irWaMEVRBJOUs3fuJjH64LJpGBlHKWQrJ3Dx7+bMTQT0PrXd2altkidtxKzecYLc0FVWu7YQ/qjFKWULxOUG72i+WlViXr9Ci0IZIAO90iGQ8qTE1bTGfl0znw+Zzabcpat+TDPSa/W9K4yBk5wFAQcphEHQcBIKwahYhQFDENNGkhC6ZUOVXu/rJCUDrLKsspKFmXJoiqZFSWXRcVFWXG2LpkYwVwolkKwDiKKsA9Jgh4N6B2MSA72iZIUGUQIqXDSgTBt6mCTXrkRoR2l3YIxlmyxZnwx5dnTC9bTlccseOmW3Fp8W46v9g3nk/5SazkwFV8NBd/rRXwjDRmV6xrvv2rnA+GVX4XzZX9JWHPSpsywayFLECHGBcxWJT96esZVKfhgtMe7/R6HzhBgqICV0pw7wWfrgk+Wa85FyFppRD8lOD5EDvuUgcJIt1kDN/CtZv5ep4rJgu9WqDVWiho11daIqTUP/VJ6QL8YeYyE3X19qx8A4G3uBXAbvcIS7OyhBo+8ff9VUMAdN6zYuc5Nm6W10+ruYZvPHR0xdfOti9s+uPbhm0Pd29pywb/eLn9d6+Lln1tcm4mxUQScq6vUlIRAUYaK5GhEcHJAPp5Q5iXT0PKbcsUPx3MO05BvDkOEKRC2RCnJnWGPD05P+fGj3/LzZ2eoMODh4QBNCUWnznl3JI0Q74YzqMAJIiW4Nwj5m2LAtJqSLQyVKTjHUUjAaa7FBa/NQNeiqkWdkRSLkvPqgvV6zZ2TA/YP9wnjYJMXsOtyFM0M+hJCp4RvL6w1Lgrp9SKSowNsXlIu59jFgvV0znyxRmQVKs+JnKG3KuiRETtLgKWnJIkQxAJCfFxb4RPCHAojJIW1ZM6wcpYcQe4kKxRLJVmGKYUOsXGMTBLiUY9e6kMVOk0QUYgMFU6pegyN1b7d4Ktbn97Y/9ZYyqxkOp5zeTZmOl6QLzOckWyeWXd+xeaZdvgBuBuWu0W7ir6p2C892t/3R33+rB9wtyrpVRWhtWjXEaiN8NcCEWmf/U8N+LP1uGvAoyBkvDJ8eHbF59mYNOhz2htwHGl6pkBjyZRipkOerAy/ma44MzCPJVWiiA9HjO6fIALlhXQTytjhZ8393VCncp0ajwq+M6XQGivlxgvoXmUMvF3UhkFEZ05eXVYunBPd5f3G0b+CAuA3q4Ptpn87n281VGgbyr7uXG4z8s2ZvQW2ey4BbVOb3dvYPetLHIn8KaJjbUp9Xo2RANs9cF6G2/ByEi0vbtZBA4jjHDgpcIHCBAp6IfHxPtX5PvnVjHmheVxpfjpb8dV+xNeGhwRaQ1UhrGEURXx1f4+LsyGP1wsGiyX9YY87QQw1JsGm7K1zP/VsbAMG1TFeZ4mV45v9kHmesrRrlsuSvLLMNJQSXIszL+o6LEHbIeTaYqmVACdxBsp1xczMMHlJkRtG+wPSQQ8VBiAtsoOn03hrrOjYdzXUlnACrQIIQ0QSE/VD2BuSH6yoVgVVlmPWa/IsoypKZmWFqwqoCrQV6KpCGdNauv6Sdbi+PwAAIABJREFUdbczAU5I3zAokF6Q6wCnQ1wSIeOYKI6QUYROYpJegtQKGSiEVjgl2mnZOErc1uyDD3tsoiWOqjKsVxnTqzlXZ2MWkyVFVm2aSdTrZiPsGwWr8wy6Mf+Oh95n8Dtia9izJe8Ky/eHI77Ti3igLCNTkBhH4Bqfpb9D6RrDXvvEP+HAVV0XDW3yoQrIkbxYr/hoPKGyBQ/7fY7jkAGW0FZIoNIBF1bwSVbxSV4xlQG50thhH31nn2h/RKWaGL0fdzeNpfZZ3VzcfIvXUuD7JkgV+h4aUtVP3D8keftX316yrqPsN1p55/UWvfly4I+sADSufNeiTG1Z3I0VJqgnuhbVzifSbLD8PSN8uTt+w8gbIUPjE3C0jH5zFxsFYMswbk5Vk2yPftU4/wSoA5Byk8167fCOwvSFL9kRK503N8+j7mrmtMLFAWUcEB7ukdw9Ij+/ZJUXXJiI3+Q5v5iu+O5+j3f7kS/FcZZYWO6mEX9+55T/9PwRvxtP2EsSDu+MkDICl7Pbp2BzEze49pzFYwNUHEch39+PyRws7ZpiWfLESqZWUDSK/q0K/64C2wgJrwWbomJ2taSsLOtlxuigoD8aEKUhMpR17prfEw6uoWs1XjIBSOGtU60jRBQS9mJsZTCVwRQFVV5gi4qqqqjKElNWlMZRlh7G2ZmmzW9DEmqkOKkDpNZIpdChQkcaFYaoKIQgQAS+qYzWAc2etk1IRLC1ZzdW//ZvcFgLRVawWiyZXk6ZXcxZzlfYwtU8oGv9d+bUdRSxrQs1ioVon3/T4W/PlLwjLN/vR/zVMOH9EA5MQWpM3ZVv42UQOKT7/9l78+c4jizP8/PcPa48cZEEb1JSVUmq6pnuaZvZMWvbf3p/XrM1G+vpqememS5JJakkVZVuHgBBAHlnRLj7/uARkZGJBEndVIlPRgEZiIzDj3d83+UgMiHtL1ZB+DdaSzWvEoS/NwkPx0s+Oj3ji/mEnSjl3rDLQSRkLkd7R6kUMxXx1dTy8SznSyeMogibGJKr+6TX9pFeimuVMfBU+mXFI79Bv9VqhMOVPILWCTpKkKp6pvcrEwnP35jb83ugeh2tGRA/zzH6CV0Amwy4DXW2igc3hy9WVm63mN1+j9anmoGy6RioT3DfwxRuRx5eUU1tIdsqerMRleyUB2NQWUwZLYj7HdJrB6Q3z5mdjzl38MBa3p0ueO34KQf9G2Q6QZcFuJJMK964vs97k3O+Go/49PEx9zsZe92Ui4WBWGn00vyPtTn0ZcUIFTdSwz/uZiwRSjvG5wXWKsYoCl0x/jatQdAt9bHhGWr1z1vmowXLecF0Mmdnb8bOwQ69QQeTaFTUGrO169b3qmrRt9Gc6p2UjpA0wviUxAb1yzmL9R5nJSAjpcNZWykAIKptrkuoFqcNohVKJFQRjkKDLldD0tVX1iBTqVL3qnRMaWa/VrIqpd57sB5rHbPpktHpiLOnp5ydjvDzKk3R11HF9T+3pshut4Ev8hrlHWlZsGuX3BbL7zox/9fegDdix4EvSF2OCSFx1ZUDEqTEhbziNA7Qf5Nm6llBmipY02nG1Gk+Ojnm/ZMT5kp4s7/PrThiF0fkLVY8M51w7DSfTGd8uig41ppprPE7XbrXD0gPdrCtyH+p3RGy/qbfiOtUYIhXgo4jdBSt1u6a7vSKl8GKR62kRLXLGlfMz1MJ+MmbAbWHLNSfr4P9toWwSIUewJY4vtYF26Z8c/G13h8rwGzFkGuI8tsZ8D/PBfDjUT02tYdy+yDXAkQbQ9zrsjydUsaabH/I8M51Zg8eU7gRp+WSP80X/POTJW9dPeT1LCVTIG4J5ESdhLcPrzJxBV9Oznn30RH/9Jv7GFtWaYHtDm2b8yasqtzVLoMS8QuUTrjVjfi/JUHZgsXRjLIsEK8ZS0wuijV7bGsRlUpJbAsuqSrSOYXLHZOnI+aTCefnI65c22OwOyDrpaE0rqZJnRV807FxXb9q2e9K4WrMRVajL0YHBtCkdtRsTNbcYVvLQnvwPtSBFJGgv0izmxqEp/6uQLCcUa3nDcLaV7lntrTk85LxeMzR0RPGTyeU87wqa2yqG7Tz+m3rnVfo4EVauXTwoJt0v5xbPufvewn/da/Pm5mwX8xJbY7G4sXhNYgLbhGFDRkZaQrVPDRv3IYNRfBRjE97fP71ER+fnfFkadlJh7y+t8M+BaktEe9ZKsO5yfhkNOfj6YIvneUs1ZSxJ7mxT3JtD91NydXKtNjGZV7I71/PHWEoXTVvJjboqteC/dZuvV8G+aYWBo2b7OfM939CBWDFJmTj6Ko6Wc2YBPG17/6bXH+zOKXHr1jhii20b3XhGhev+oq+H2rcABuLwAuhX0Cny8IYCg1RplH7vdAueFmwXCw5KTM+WVr+25dHHNy9SWJiFCW4AuU893f7nI0HfDCb88n5Kdee7HKvn5BGMWI9oYMerAeW1hBx/bGSMK4qluNyjIL9RPFfdlLOnUJOc/Sy4EGhGHvIVQWgy4WVvUIZGj91W2iplWbrNbYomZ6OKJYLzs7OGOz26e8MyLodTKTQuu4q2Bgiq3s0bg5/UQlZ+7juiql3pZcq+luqeWqjbbLal7XVL63vti+9+Tn89IGROqkKL1qWi5zpaMrZ6RnnoxH5bIktBGxVQreZl413qYX/ZTHva1UOHdo5Os7SLwtuUvDbXso/7Hb5dWYYlgsyWxC17Lw6RVBhg76SGuhEVbOfKvCvgYR1UGpMRGkSRnPLO48e83A6o5N2uLu7yxWt6LsSYz2lCBMivvaad05HfL4sGJuIIjaw02Vw6xrxsIc1gtVV6t/GXH4b0eOoFQBQkUElMd6oShVeH+MVXvfLpjaitX5crRTonyH9BAqAu2C+bxezVVqYr72RUvG0Wg14nije5mLY3ECranVeVUFKVD6/tTldffi51Lv+OZBUEO5KDWxZUFoTZ11UkmDNgsI4okGPwb2bnJ9NWC6WnDrHp0XO/3g65c3hFLOTsR9HSJkjtqBnEn5zsMMiz/njyQl/+PIBu/duEHVjjPFgXfjXVApULeFWr5VKSNfLx1vwBZlobmaKf9pJMFaIRjmyWPLQe8bGsFQmNA+q3nTNQl+z/GFlQVbPUJMD50sW4znFImcxWTA+ndEd9ukPe2RZHKw3o6qSwm3ItkI46hLO0tyRusWpr6HrLTtKmv9Vf5Eaal89n6xB70JdJKoB4eqaCjUK4FVQLix4a3GFYzEvmJ6PmYymTEZT5rMZeWmhrMeiDelvPGFT27+tALR3qG+eIaQ1OlJfsOsKbvmC3/VS/nGY8mamueryEPHvQ3PE+o7K+1D9TxySqCD8Y0/oetjuj1BpQVrjTczEwu8fHvHhaAYScbPT5143Y8eXpDYUpCok4kQMH47nfLwoeIQwMwaymPjWNeKrO9CLKHWNTn57QbNZzMcTrmmyBJVGeKOa+Jv65V114oukE/5SqA6KhZAeq9aU3J+fIvBypAFus5Sav9FYJuum4nb//7OnokYWfMg3d8Gn4wg+zC3o6Sv6gSjUIl9Bs3Vp1UakKEWSZOgkpdBTClWiU0Pn6j75rWtMJzNmecFjFH9azPn90VN60R5ZnNBVGmyBkiVX+in3r+7z9XzJF2cn/PUoJT7cZ7cbIdjQVbC95C40y6mVgBrq9Ygt0OJITcTrmYFhXIFWOTpf8tA6zrxnWXcQrN5xJfBhVSuA1t8376sCUuDBLi2zfM5iWjI7XzAdTMl6CVk3pdNJSToJJjYYpUNlOtq54tLoH6uyzawSFNYeTdaepS50eOkcNhX61l9BPE2yRX0jbx22KFksCxbznOWkZDaeMz2fsZgtQmEk70LhnDXB34hjVk2J6s9snNsaTx9QQPFChCV1Jbsu545y/F2a8I+7HX6TKm5Q0s9zIh8YoiAB6ncejUPjkBhINSQAdTZJ6/EEUAH6nznhy7Mx//zga85LuN8bcLfX5Zr2dIoC7YWFMpyL5sul5Z3Tc770nrPIkGcxandA/7WbqJ0OZaSwmiYAdHN+nkXPOsvhsUCaxKg4Aq1war0C61a96xdOvulpUn3+mcuKH14BcJveennmglqtuVrYb0L/vmJWl4/8NiVAqv9qY8sLOMUqG6HGUn+GWtzPmYK1uD7mHkJ/8jjCJDG51pRKsJEi6sb0bl+jPDtnOpsx8UselCX/cjZmrxOx3zG8nnXATcFZVOQ4GPZ4+/oh//aXcz54dEQnTYmTvVBK2FbMvDZ3nsftWpXexGs6xvFaRxBilFbEowXRokCs50w8C6VDB8GtnKKFfLS3SfNrja3XQYKCy2Gez5mPJ+jEkHYTuv0O3WGPTrdDmiZEsQ6ogJEmtKDeMRfUjLq2fuuW27tvbj5//b3gA6gtzCZj0YF3grOuqh5YUsyXzGczJpM5k9Gc+XhBvnBNBp1vEJhNgd7WLOqHfJbyVB9zCBbjhZ4t2PdL7ijP77op/7jT49eJ5qpb0i+XJFgUOnCJajyUd6F+hAHSCBLDhWZKNUqhAB1RqpijyZJ3Hj7iy+kp17Lr3BgMuZ4lDFxBbB1WRYxNwtel54PJhI+mc44izTzRyE6H9NZVBodXKJKIUnzlkPjmfGnFB7djrA6HTiK0CZ0pA5r9iv89k5qpWO0mv4bgrU4UBCWKlyDU7lL6EZ7M4tfwp3UY8dnk15iRr+J8nquQXrBaPLg6jkAhvvJ2SbA52zEBr5b/j0dt+863/wlYBGMUURqjIsEqRwmUkSK6NiSaXEPNptj5Y07jmD+5gsHphCtpxO1bB8SRh3KJuILd2PD2wR75yTX+5eyId5+eY5KMt64M0CpU/ENqJKBu5KJXi6iGRX39tJVQtg7RBd3Y8LooOiphN4mJnoxQ8yViLaeSMKfuIFiRp9oCHrDrkNNmKdnatwyrKNUqQdsuHdPlhOnpGKITsm7GYNij1+/Q6aVk3RQTacSo0O1NqnTCWon2Aq71KNDqjtuqaeG3CeUar6n2lbcrkMQ5SuexhWOxKJhOZ4zHYyZnY6ajMWVegpWAbkgEmFaq/jPQwDVFYIvF3zDiIN6Ut2jv6PiCA1/wurL8Q7/DfznY4b7y7NqCji2IQ1HncNna5+89Bg9ioZtBkgQlzdnqmev7CKBBKdAxoxw+fjrmneNTeirj9f09bnZThhKgf6U1YxPzUAwfLhe8O5pybAzTWFN2DN3DXXbu3YRujDOqqpZ4yXA8h1nVeynA+Csh5Su00wFxmqAiE6ajdtVUPzfdBr9kqsdEiazxA8FeYoyu3Fe/6EqAVXHMLSvpRbRa2Tq464htC+bcdkJ9la23EuoQn1dL/YemFxxhIViUBAYVpQk6jrESWkOX2qNiRe/wADmfc/ZkRF6UPI0SPspzfv90zK0s5R+uDDEIUuaQWzrK8Ns7t/k8X3I6mfCXoyP2IsO1nS4KhfglTT53XanvubLIBUGmLXEkXHWe/+g9+dU+8dmUeLzks9zy1MQsJaLQmqZgUBumWrt2daDhGVviu0MPUlbKiIcSFuMF5XzJ2ckpJlZEqSHLMpJuRpqmxHFCFBm0NmgTmJkSQUStCjy54Aeu3QZrZXkFvPONjPU+7BvlHGVRUBQFeZ6zXCxZzOYs5kuWi4J8GWoP2MJiS6iB9mcG7zWDfMl8bDu1/sVbjHckztKxS/Zswa8yxT/0+/x9v8Md8ezlC7quJKIMqX0EZh7krUOJDY/Z6YR8f2EL6lC9g9IQJ+S554MHR/yfR8cUxvDmziH3Oxn73pHakEEw05qnEvHJdMH7owlfWs8ojiiVEF3ZJ7l1Db3fpdBSCeXVezfxoc8YhuePT1AAHeCUoOMETKjO2IS9+I0vvKLnkKyvzY1EoJeZfhxs4gU0ye1nbIOuVnb6ZRrq5XziokLhWS958op+SHo2xL6ancCgShwqiZogJest3oV2s1G/Q3bjCvnZlOnyUybe8NDCuxPLlUdjjEl5I1F0Co9xc3QEO90uv7txkz9+/YDHownv6Cf8fdphP06IlEdc/WyV+tEWKs2PiiPL6m/iHVpZOhFc957/pCEZaHqi6U2W/LkoeaozRhKvMgSsahXz8S2HfB1V3Maj6nu2cJJaMngV8HbnQlXB3IGULJVDDMziBToaE8UxJoowURSUAKMwWqN1KNoTGYPSQfCLktCPQFwozVu5CTzgytAQyJaWsixxNtw3z3OKSgko85JiWVDmFus83lV++7oz2EYg7voS8Zf8TVqC6ZI15GvhX9KxJUOXc+BzfpNq/n6ny9vdhLvas2cXdKv6/krqgsOeOq1SUSKRQBaFqH8Nq/oRGxqbDqV+rcS89+Qxfzg55nGec7W/w2/39zhUnl0bygkXyjDSKZ/mjj+O53w0z3mkDBOj8f0O2c3rJNev4DsJhQanfEAAoNU99cUFs2oPp9Qht8Er65WgkgidpYgx1NUkVbX2XgU7X05tyF9aaYE/R/rBFQCxF6KdttOaBl+pvgI0PdHaxVu2jHh1+JlzUZVmlWfCjK/oJ6EN68bjseIxSYJKE4gifFlixQcBZTRmf0jv/k2mp+eUdsSo9Px1sSQ7WyLqFHfQ5yaOnbIk0VMkE+4O+ozn+/zp5IQPTs9QcZf/fLjLMIpRGsQWhBD0tsnUerjG/8fKXPIO8aBVqA9zC0fSEboqoqc92aTgr0XJAwtjB0sRrLRSBdv+/3Y16YY2heTGsbptbxPHoKAq6JMvSxDLXOWgFUoptBKUVmilQvMho4miCKVVaGGqQtEflA/td51venJ4G/L1bVmGn9binacsLNa50JzH0yqHXLswWq4Mali74aKXUMv8bd7Zs5lFVEcgKu+JnKVjc/Z8wS0NryUJ/9jPeKsXc108O+WCzJYY74LbghpB9CgvQSGIQFId/P7a00T7t1GA6r28jlh4w1dnC/7t8RO+nM3ppn3u7+xzO9YM8wWxs1gUUxXzAM0fx2M+nC/50glnaUKeKrq3b9C9dYjZ6VNUbXmbwj/VAIS8qBePyV+N3rqb0wtgNHGviyRxaAbUus8aOvWKgJWxuRJmq66Qz/JUvez0ckUnVJtcXGt4JfQo9+Lw3tKOWHrRugDtSdueyBc2uH+FBfzAdAHvvvw8AURQcYxOO6goxi8WTfSyiGDSmOjaHunrd1hOP2WRlxyXlg/LEvtkRGyE/9CNeB3NlcUSk58SZwNuDAacOs+jh4/53199xRWj+NWVHbpRVvnFWwpnW/A0j7eB33uom9uIVqSx5ro4YtF0dEY/ihiOLJ1Fwdel51RgZoTSSVPedUUtBfdFhqtJwG9biL51vOVOcCHwy22zolWtPVf7S4IC0HRoapQg1QjcZivVyAXCqoDXtq6LbWSjxpu/DW36T4K/P3aWYVlw1ZXcjeDNXsrvhj1+nVbBfsWSxJVEzlaBflULYoITUCFILEgnDpa/ohL+1YvWypqn8vknFCQcTwv+5YvHfDpekOgO9/v73O/36JZzYlfiUcx0xGPR/HFe8G/nE/5awmkcsUwj1F6HnV/dIbqySx6HgNc1Hue3vPt3YFQeQZmIdDiEOMLXSFSF9rzigc+isCfabdHXf6l/Xx2QZ/dB/0npp1AAtprwDdjp61Sf+vg2uH8THq2PPeOm4tcSiJrvSN2bIBT18Nvbabyi70zP8GkDa5YHwWZBwGvQWYJJEopRBUX7YB1ZI+heyv7rt3jyZEReLJmWBY/E4/KC3tkEiXZI+h2MQK9cUk6n9LIuNzsDHg0tf376Jf/z60fEUcQbB0NSE0ORb8DwtYfcNY8alAC72uy1ouCCEmDQXPWWrvYMehHXTMrV85x3Jzl/sTOeFJaZTlh6g1WVYNlcds3SfkHFqUEn6n8tQe9ldU5dbdO33A11EF/7VuVKMITvtvZafW7TYlNffE5pn1sL/c2Xew7VvodG5tcfHHgd/PXektqSQVlyy855M0v4j8MOb/UzbsWKoc3plgVpFRtQry1c3R7MBUaoBboJZLpyq2wWipKV20YZrEl4OoX3Hz7l3SdPiFWX13cOeGtnyFVbklqwoliYiCcYPl46/uVkzIel55EyzGINOwmdN+8RHe7iujG2VYRAbQj/7xqg3wyjKIgiokEPolUA5ssrpl4eatfUCKunrhi6SY7AHyxVUYuXkn5wBeCbitP2UAo1ar+GhXGJDvEt6ZWwfznoolvGewm1ypMIlSWgVOVPDj25rQciiDope2/c4rwomOcF89GMJ87wYZ4TjyZ0lJB1MgQhsQ6VF/SU4d5wQJ5f43h+yv959BDrLG9f2yVK0iD83Ea+d/1oz1oylV6AUkgCmbLcn5dkqWFguuxnCbujBR/Nco4Lx7mOmGkdYgMUrClIth6XWgBvCmJWn7fFw9QRy2EwW9+r2yK3LfQNYb/2+zOU7XaAcy0kv/fo8bYGUPviXSjsY0u6tmTPWa5r+F1/wN8NO7yRGK6LY1gsSJ0j9i50Oawh/+q6ynuUeIg0ZAnEVfaHr5i3qxl+laKoNCiNUxlHk5L3Hp/w7vERqcq4f/WQu70O+3iyIuQ2LpThWCX8eVny76cj/jTLOYoT5pHGDTKSG1e58sZd/KCDNQpRslJQNkk2DaEXREDb5X8BpxQqiYm7PZyJ8FK3Ad5yvVdKwRqJBN5Tp79WR7dqZ5fhzS8T/cAKwAlwANsTi59BbathA+pvq6nCd2Q29SS2ru9Xj/uqC9aPTC1LpOrbFID1JEJnMUQaawsg1KpX1b5zsSK9soOdX8Mu5izzgqm1PC41H89zdvSMXdMnNil7FBjn6TnHDaPxOzt87EseL6a8f3JMEiveuDJA60pYtP3/bcv6AiOu/lVrUvChG6wROqnmsHBEODqZZkdlHJglnyxKviiXPLGKEZolOkR+14GAtQVdX/fCeLWE7WVrtT6nKePbeuTNAgAXvlu7QTai9RulYtv3vgu0v3mpWvDXzxn6Mihs6ORnbRD8WO6nhje6GW/3Uu5EiitY+q4kcZbIOVRd8bBBKULjJKVB4igE/Jm6OthlAljwKsJHHZ5MLe8dn/HuyTkjFPd3Dnij3+Oq9qSuQOGxCBMxfL60vDde8sE05zGKuTHYXkJ8uEfv3g1kp0seCaWueM+mfkf96BVy47aN+2VD6Jufdf1/Hyl0EqPjGKdr4b/lnpcMwy+RmtTIBg1sNZWXCrFsu2d+JorTDx8EuAqt3kLb/9RuC1ovwVoo1NPgN6yTF1+oNfMK0ye+LvzRlAp6Rd+Etk3htxjEze6P9SZygEQanSaoLMYuF1X5zZWGbY0QDRLSG/uU8wXFdEFZlpyL8HWR88FkwUA0nb0hWgk7viBxnl1KVDdlyQGfnTq+mk3xjx4RRZob/Sj0DBCgrGJPVthfSzhvvkB13AXXkghIJHQFzLKgY4RdpbhiYm7kER/Ocv6yKPnalZyVhoXSlGKworCeqjRrW0ndtMqfN/abkPzlX13/Y62FtY97WvzvkufZohBcOG9z0bQV8A24pVICpGrGY3xJ7Eo6vmTfOu4lht8kKW91Yu6mMTeNZ+hCK1/jfdXEp8r1aZodhZWjYkHiOBT4iarcLV91HazHvK7ApxTeJJQqYZJHvH90wrvHJxznjsPBHr/e3eWGUXRsjvKWQoSFMTywwh8nc94ZL/jUKc7jmCKNiK7t0bl7ne6tK+SxolRyQa5LG71pj7m0rc/nUzuAzUlQeKJOhjTW/8WZuwQP+MVTGz9araVnnf1yawI/Uh2ATTN9U7O/bKmtjquWiFZtRnzx1GdQO+VPoGow1FRsb/OqV6v/p6NqTdQgkGhNlCZEWUp+PkLXgViVVWMFciNEuz2yW4csZznT+ZLFaMG5Fz7Lc6KzKb04JeklaGXo+yJ0hMNyd9BDnOez82M+Hp9jv3D8053r3BimZFEMvgCKFSO+4BNgtXi850JdelFIokkoMYuc1MMgTbnSTTnMIg4nCz6ZzvliueRpqZgozUwZFqIoxLSYziaLZou1vYXpXDjlBRe3r1OcWj0NqnFfD4T8pvScjbtmAHjEWyJvSVxJzxbsSMmhgrtZxFvDDm92U24bYVDm9PKCxFuiNp8gPK6qkBmtfPC0ZFHI8deqmuN2bf/6vR2IBpNSqozzQvH+0Qn/88FDnhaWq4N9frN3hZuRplcu0K6kUMJUG450wvujMe+OZ/ylcBxHCfMkQvb6dF67TufeIfQ7FKrVifRZo7WhS31ThLJWAKIkJun38ErhKp74it29GAm+BZytZ1c0tJowL/KdIOofnH54BCDkELUGYTMUr27L29qstQDYuim2LdgXxVy2TNaFU2qocNu9X9Hl1Gqt/F2omnvXwNZqpQB0O6E6WhEq7OumYlkVr6Y18cEOewiL+QL7l6+Ze8+xB4oSdXRGT/aIOgbRhj45mSs5EEj6HRJ9lT8+gT+cPUZLyX9VN7kz7BJFvvIHt3P06vdsBwbWArMaB9/i2K5EYoPWiu5iSbqYkbmS/SzjbtrlN92I95+O+WSS88CVPPGWcxUxFaHANz0FVqPbFlL189QKh6/g+0sGuOlE+LyJaMUKSBX9386FVyEQb2W6bmDGNadsFLYWilAHUPqNoNC6eQ+eUA/SEXlLryzZtSXXpeSeUfx22OG3O11uxppduyQtcowtiTZh60Y/8yhvQ4GfiBDsl1QBXL4I7yWu5emoxlULqAirMkaF5sOjM/6fT/7CUoT7w11+Nxxy10C/mBE5hxVYasMTlfLe3PI/nk74pHAcRxHTREM3Ib13nez2NdRen/lm24N69LcJ90vaHbfZ67bv1X03POC0oDsJca8T1lUNdNQK99Y7vKKa1kvG1fuu/tn6W1jv4tzL7Uf+QRUArXVI3PvGMkGoU1Ig1BlvWKn3TcnK1WXbwMwzrlmfugYFbty2Okc2Id5XW+M59D0pus1lBF9Vu3MoVBwRdTNM1e1v835OwCqhiBXRbp9rb73Ok9JTfP2E6ekE74SoKPjXJ2fI/oCyG3FLGfrwKNZGAAAgAElEQVQ2Jy5KespzvZNQHF5DH8Pn41P4/AsWh1f41X4VGFjkSGlZj3ZvC7AWGtDwhSDImnQyrZEsQhvHcFkSLUekohhEMVevDrk/tPx1XvDpLOeL5YKnecFMKZZKs1SKAkWpVEjl82bDd7IB9z93Sp4BxT/v1Au0oXBsIv81ckD9cwNN8cG/L4CxlshZEm9JvaOPYx/HG/0Ov+7F3E01d2PFoXf0Fksyl1epfa5BLWoTQXnQYsN+N4RCDZmpOF+lpDXITj0EtQsglPi1OuXx1PLe0RH/9vAhVjR3dw741c6Am4mhb5cYbymVYqJDmd8/zhb8f1+f8JFzPIpjZmkEgw7m7m1237iN2utjTf24snH/7cP9IiV6L/9LcDHoJMN0ukgUh+tVZW2dX6nw27/9iuAC10FEVevWXTgv9KLyL3MSwI+VBih+5UPdNOtb6m9LWVq1paytdo94QXuFFwk9hja15mc/QfD313f0oYJbnQbY3F+kyQ1uYRLf+I1/efT9KABrCHsVcetFQBt0lhF1usjSQZmz8hEAXnDKU3pBJYbk2i478zuMPCyKkrmbc+I9H+QlajyllC6mE6M1dEtL4h17PpQZjvZ2+Pik4MF0Co+eUFh4+9pVjALRBdiCCylvsA6NN56mtvVbI+oq5JsrQzcviYuSrnf0JWY/Mdw2CW+kMV8scj6bLniUF5zYgjOnmCrDzEcsxOOkzr3Xq4Gr90yTqNxGs1rrWDZ+rjTsZuwvTMoFV8IlIkPcurXaFrA1U2wqH1b1E3xI50uspeNKBtayi+VACzeziNc6Pe52Yq4nsC+OoS/olCWxs0S+ruVf8Za6nn/9TxwkGklMiPY3HmRVBKjSGJrvhssEn7/TMQ8nS/790RPee/KUsRVe39nl/rDPrcQw9CHDwIowMREPRPPevOD3T6d8UDgeRRETY7C9jOjmATu/uYW5MsAmGqfa3LDdHZOmO6nyoXDZmvPnOUalq6ZceVqtn8OURJ0U08nA6PXryCUR634t/PMVIa09XhdVhjUErvpYt7L/RfcCcLYy5psjNSZY7bq28r0ZqcwKgQxfkBVD0y37fcP42SSpvlsrACvr31eaW90NYMW8ayVg/Srfkraq89/+ci8V/cDvEWbF45VCxQlJr0c+nuKX1ZrYqNDlFRRGEInIru9jlzlumVOUx4yd4yuvUPMCxZSOgOkmXFcFHWdJrGNPOSSLWezs8eVIeDyf4R4/IcZwd9gni5LQVMfmK8HWtAj1qydZi5Svx6nFJIQQ3Kg0SjymsER2Qc9H7OuYQ625EyXcNoov8pIHRcGDouS4LDj1lpHX5OKwymBFVw1e2rUuGlV38yFWtIZybSo0vnX+lu97Wb1vg3i0jm0TJ3XfDu9QPkTmB2U8NO1JnaXvLXsC11PNrTjiZqy5nUbcTWL2tadPQWoLIusxzlWdFWpEoQoWlFoBqDoLxya08jX189nVnNXCv2Y0KJAIr2Jyb3gyzfng6IQPT844L4VrwwN+M+xzGBt2vCdxHiehve9j0fxpWfC/R3Pen+c8imImsaHopcRXdujfvUHn2h5FaiiVbyr9rVQAaYa2rS89b4u1BXmbFYbv+mY2nFIkWYrJMrzWYR03+unqTmv3eyEk6WdGLwx8bTlRaK1zGpRy7XxZNx9fZvpxugE2fbzbHpRaFD9ndUkFk0m9mF9kS2y/UKMESCvm3yvES4gU9q65vmx89xX9WOQv/BoYlAQFYNAlP4lw8yXKrm+z2tC2WigQTD8ju30Nbx2jZcGiPA6XXC7x0xnKWUTvo+KYQ0o6Niexnj08r/UHRErzxfkJX0/OWcw+x926w82DHXppEoLGyyplbC1VsE3V+pbNNVufaBETkAAxQm9hycqcri0ZYNg3EYfDhPs+5VFR8OVsyZezJQ9zy3HpGDnLxCoWSrEUjVVQKE0pgq0r8Ul7j11E2i4+02Vrfds+rRWAFoq20p63DINH4zAulOyNvSXGk7qSjjh2NFyLNNeTmHudlNtZzLVIsy+Ofl6QFjkxBbqKH9CV3R8qeHoEi6IMgl8LYnSI8I918OU3hVku4yEKVAw6ZeE1j6cL3nt0xJ9OnjLxipuDfV7fO+BO7OmXQQnxIsy04YmJ+XBW8G9nE94Z53whhlGSYDsafbhL9/4NBrevU2YRpWZVAVJYs/wbEVwrS5fMxjOpkUNhbXrAKhWi/7tddJpWKEHV/aA1HFuat/+C6TIDsKXoX0Cz1/7ut++bl4d+eAXAAb6Upu2pBGb+7fpOV8z0W3w3RAGH0t5B9VBVG9MVCAe1zbR+7PuiumbUy14c4ienFhBUM0Qngoo0ybDHstOhmC5xrqAdZOsrGNd7RamASBHvdOnfu454z9P5lOXZnDPncLmnmOUUT86Ir+yjooSrXug6T8dZrvicNE3oyAF/1RFfnR3x/37+Nf9gHW8d7rKfRmhxUNTZAb71xGqDN2wwgTYi6MJ6ltiANpjCohcFcT4nXeR0TcSBMdxLDW+nHU4GGV/PSz6fFny9LHic5xyXjnMUS6OYY5iJYekdVqri1t4HJVxkvWLwNuiszcOa8r6WVfdBvfHd0LaphvIhWJW1YiRqNYuJt8TO0fGOri3p+ZKhCPtacS0x3OrE3OlmHGYJu2LpOUvmchLnMLbEeIuIWy/D6itBJxbEYepGPmlS1fJXldBfIS+riWlJYdGBr5iEwsc8GC3416+Pef/pMUal3Nvf5/XdHQ4jzU6Zo6uuiAutOdYRH5aWf356zvuznC9EcRYbylSQ/T47r9+md/8GbphiI5rWDa0F0fo9cJ9vy5jb3/VV0KqT0EAr6feIe92m/a+7wOKqcsjf8t4/L9pEt7bRdgXAN43C2nKi+r2Jq6j2hnj/iy0FfHIC/R2HfUGJ5/1mo57vk2rgP6z8y9yXPyS9tKvgJaP1cZKGaXsRdJwSd7vY8wl2mV8AuesreAmZAWIUZtihc/cqxXLB9MPPyRlzrgRfOtR8QXp0SjHs85vMcMPE9H1O7HIGXuGSFG0yEtPlq7Nj/v3hQyaLKX93eMDhMMPEGlUsL9YKeJZfSvx6Mkztd1YKEgUmwiwValmSlAvsEpalZkdHHKiIax3N/Szj2Hke5yUPl0uOl0ueFpbTMuc8z5kiLMVQeEUpQq4UhYRCQ84rRIJS5SoM2NW5721YugE2qlgZpLIQQ0CjNC40i8IGSN95IsA4hziLFjAiGCBzjoES9rXmahJzJe5ytROzF2n2DewrGOAY2AWpDQiBwQao31dFeip72VdR/SFE1IbUPiMQJ5BEwdcvDnxd1rk14NJyj4gCZfAqwqmYYgEfHT3l3ZNjvpjP6Ogedw6ucKff5ZoS+sUSbR1OKSbG8FiEP81L/tvJGe/Pcx4qwySOKBOD2u0y/PVdsltX8P2MQssWodtaFt+Y921bX7V2FNaiI7goMJruzpA4y1a1/zcu9csQ/G365hzZr+3xunKMgOiVZdre+i+5tfejBAG2XFptG+kb03cJpfCVxlt3/q6VAS8/nsb7kq+Fl4Nku+hUBEsGbYh7XRZJjJtOcWuozgrHrCufFRq8KMxuj/4bt6C0zD59QHEyYjwv+dp5zHxJAczo4HoxN5Sj50oiHENn0SoiHuwQCTw8P+Hj0xFntuSNxR5v7ffomRRRRcgQcO2goIvvVvuqV+e0ha4DUcGC1RplBJWX6MJibElaejJxdMSwp+FQC/czxSjJOLcpo7LkaVHwZGk5KxxnpeWsKJk6YeqFGYo5sAQQjVMK5wWLxzXBtUG0h5BwWz3lakbElSGwzociR0pKNCXKF2gPifd0gK6DBEemoGs0vUiza1L2TcyVSLNnNEOlGEZCKpDiyXAkzpI4h3YWjavuBeIsdaR1GL5Q6EeUhyggKBIZMCZY/fU41yBFuyxyMx8KVIJXCUsizhaeD7865pOzp5zmOYOoz93BkMN+yp72dFyB9g4riqlJeIDm/fmSfz0b8+7M8pVEjI2myCL0/pD+r+/Ru3cdtdunjBVWBev/oqeoxYO+oRLQjEnNWTfcL55QTltlMVEvQ0WGskJhaX+zbgL0i9ECXkT4X6h6haBYc/l5D77u7Kl8c5xaWXi56YdXAGxYgwExaVlHwUHVGtk6quIyq0kuzNm30ZdX5ZvlOykU34h+MZvq+yFhQ9nzLWVNKeJOB93JcOMxrrDoLf7SOvfZAaX2EGvivSH9+zfBOWYi5EfnnHv4PC9xyxw39hjl8L2IGyaiX7WN7XmL1gb6Q0Tgq8k5n40XjPIjpCy4v9tnmMREBqQsCUVloC5du3opuMh4/Orv9XcAlCCxBq2Q2CGFQ5UOXVoia+nakh2lyasUwUVsWESGUaw4TzznpeesLHlqPWcORk4YOxhZy9RaCg8WR2iBBQWe0jusDwrAhfqd1bMrB0YUWgQtoMURiUeLkCroimagNDui6ChP3yh6WjGMNDuRYShB8Pc8pDhiX6JdQA+0D8LeVPECgkfENzn8q7Df4ApUEUgUBR9/pAICUA/0BbdMa3VUCIDXQfjPCuHReMqfR1P+dHLKzDkGnQF3uwNe68T0xZG4HAFKERYq5jGGD+cl/2s0551pzhcSMY41RaYxewN692/Sf+0maqeLTQxOVxktzVxvKiNtiPkifSteV/8zhrjfRXUyiHSr9n9T9Jy6CsAFsPpvkXe1XUjb/9T6tHmkfcxf3kDJr/14aelHQQDc2jC0l2ag9ZKXm/7SgJjWvqnvT6taFf592Sfpl0XVFqsAtVVKpmoqoJo0I+p10eMUN56tl7SnEv4td5L3nlKBRIrs+pVgIZqIqXUsn444FYVb5pTTBYXLKfQQl8TcNIaeLTHe03E5V6MIs7NLFCd8Pjrh4fSEf/1ixnhxwOtXrnDQ69FLBOwMbA6+bGDrQC2usI1zSG25hnFABCKBxCDWI4VFLUvM0oHN8aXCAQVCoSNKpdlTmmWsWCaGmSTMlGLqhYkVJhYmhWVcFMydY2ktpXNYhNx5ls5Tel8pAe3nDWariMd4IVYKoxVag1GGRDsi5egYRU8b+jpiRwkdLWQKUhEScWR4YudJylCF0VSpf1K5E6jcc6oWSFVUv3iLtq5CWX0IpolMgPrjpBL8dRlft0JaLowtYUy1BhVRSsIo93x5OuKDh0f8eXSOxD0O+3vcGQy4kRl2yyWRLxAPudZMTMJjEv40y/n96Zh/n875QjSjJKFMNXq/R++1Wwx/cw99ZcBSQ6lC0N9m3NOzIP/t3udnnXfxLI/glCBJRLa7i6QJTuvqOaSVyer5pSb7veg4b6eLCsKFa69hAi8f/aAKgIiuAiBaBRObNKFLyG0A5R6UD+V6VcUq6uPhJt/3U7+in5Lq6dTQkptSWYEhmElFmnjQI5n0mU8XOO9Rzq19f71oSmB21sBCQXx9j2FsEKMYvf9nivMFIx/jcsVyUTB9PMIeDLGdlJuRpu9yYuvo2TxUkO0m7KZX+fLU8Mn5EUcPjvly4vhPtwy/vrpPrKrc7bJ+CVkJpTUXYnutS+tn25Il5NIqVdWsN5B6WJTI0qJKF4rgWE/kNdopYoGOEgbo0OxFIqyOsFrj45RCdSgEcm8pbRmEPp6SoACUhEDKhqotqwRiCRUYtVKVLPVEOLR4jA9C3VhPTMjPV2UQ4iiHruB44xXGC0ocuuYMNbesYhJCZo6rUgYJVQcjVil9cUSAAHwVcFiNnQeUXWcxqkZZFCiNVzFWJ5zNSv7w+Al/OD7m4XxKVye8vX+Ve/0e+8bTsXMiSrwIhdaMTMJDSXhvXvL74zP+OC/4WkeM0gibKtRej/6b9xn8+i5qt8tSewq9Xua3vS5rY2abIlDHCmzrEr2+Zjbba68kjlPgIoXqpKS7QzARts1Da19sdTOp+KxwsV7r3yrVMeCXFs589rern7LxufrkwPtn9cL56enH6QXQ7nLxDYajgcvEVx6CasO0cr/X6TnaQPsRLrgE693wSqN4WSlEtCucMkTdHlGny0Q9RdsCLyul4bIZtOIDU1Rghl0Gr98CrZl8/DnFkzGjGdhCcEWBHJ0x3eny237G7ShmVxWkzhJ7T99aRCDZ2yXu9Hnw9IxH0xn//bNPOXp6xt9d22HYi4lig3Y5lAVrtebXAolatGaRCU0ksSdYt/UaNRq6GaRAWaKKgqgIBYoiBOs81oVCQWINXgo8Gu81Ho1VilI8znucuKawlvVV0BiCeI2vrUJP1VAntNSt/eoigA1teZsgwEpR05XgVpVQDzJGEwp6WRQS5st6QhChqxr+gDiFiAsTWqE1xFlAQzSVQPehINOFgkXVMONXf1NBWXA6wqKZFvDwyYg/PHrAn6djZmK4MbzGvZ1dbiUp+1h6RY6mxKGYGc2ZivmqFD6YjPjvT8Z87uBBZBhFEbYbo/Z77L39K7LbV2CYsTSeXNHk13/TQrvar/IqnkcXUFEfxrtUgmQJ6c4QlWWUkQpxNBtj1qREN+uvol8KK3wBmbQ2xmtwowP0M4dK5HlW709HP0YdgKDP+8C8L6Etg7M65MQRMvQrzlO3S20QhZVvZqVVX36XOijBt47Xn38pa/7nRavqD3Wev05idK+D6WSUo6IR/npb57xmUgXnXbDKEo3Z7dJVNzFaM/nsAfmjU6ajGY+9RUpLPppzVjre7iX8qpNwjZKuzYm8ZYAlUYo4Sxju7/FokvB0NuHdk2Mez0fc2z/g/t6Aq1mGNgacQlxBSJmrlYBNK7t+3stssJqPVFH5RiFaQWQQq8E5vHUoW6LLElwZjnmF8zpUDhSNt3XbYd9YinUFzNX6t3ivGm+FACK2GU5fBVrig+BG6qyACqX36/7kcF3XXE8FlQSpMgrwLvj7lUCsEG1Ce14tAf0wuhL8jlURHxt4ilyiuAsgGnSENR0mVvFgNOfj46d8NR5xOl+Qxh1u9/rc6A05jCL6WDq2wGApRLHQMccq4uOl5Z3xjPfHcz4pSk7jlHESYfsp5toe/V/donvnEPoZZSQUqh60ehBeHGKv3+RZ5shlrtB6Tq2Euv9Jp0M2GIAxIeizfcV2SoKs/bigC/yt0mbhzueRb0aYlZCpFc5L0v5/sWmADUndwHXdZyIiq0ou3jfw/2q0fAXR+Erm1xu/1Q6oLcVb33vW6q0rbflqwgJbWcUDvFICXk7yzX4TRGtMp0M2HDKaTsAGQdRWtYPQWs1m0xa1UiJIDNFej76+gYo0kzhm/uVjJueOrxGWpWU6nnNelsw8vJlFHBpD3zkiX9JxlliVdNKIjhmSJAmPJiM+G005K44Yzef8atDjcJCSRAk6MogrqiqCdlUNZi0r4LKXr39pKwa1hVvh82IQ58AK2iqwDqzHlyAuVN4LAtSiXWsfOEJqmF8XOt7rZld4qRhcbSjW6AE0/vpmzH1w24lf7anV32WlKEjFGrQgosM7mKo1r1JVLduW0rM2u/WD1seENT+/ErxSeGXw1nA0yvlsPOOjs3M+HU0ovGK/u8edbofbnZgrRtNzod2wAIUYxtpwpCI+mYXqfu9OF/zVOs6SmGUSYXc6xNf36d2/Se9uJfyNtLr7rUsXWed9l891Rd8qU4qqL4YASULU7xH3e9ha+LeCqcPwhQn13jc4RX2dvynaEAltR9s3YfgrBcBD7cDyFu/sFqWsKkn5EtOP1Aug1TGtcroEMNOvSoL7lWa1PmJ+VVthbcOv9r/fMottQd58Q1a/e6nrhxGsnzXL8RW9TLS+HoI/X4nCpBnZ7pDRkyf45aLVY2bFxi4keTblpoM7wIpghl26coiYCOs9uXdMxgvsQiiKgul0wdQWLPeGzLOImypi13k6PqSsKUp0HJMmAwZJxpf+hLPFOX96/Jjx+Tm/urbHleGQYTchMxFGGXBFVUnQVo/a6uQXXvM5oyEbxzxggsWsNVA5n8uAZmgLWBXuSVC2w45z1cdwvbWGeN5U0LBrULjGh42v+nHIWjEmfCW3nQepAjdbzywSahCgCMF7ipWlL1U0f/AtsLKqNgR/u4AP0BQpksofrg1oTSGKiYXz84KPnzzlk9MzHhc5kmTc6u5xsz/gZqzZl9BmOPUeK5651pypiIde89HS8s7pmPcnOZ96OIkilkkMw4z45hV6r99kcOc6vptQVAF/m0CnVEL2h6DA+lYN03y1P6yCuNMhGgzwSYJlM+upxe/8+q/tn39TdBEQ/ObUlL+u9oEH7y3Olfimkmx18VrLfYnpR1EAGrkP1DZA/QdxrhLMYWBLCWcoZE3wq2o8FYJh1SwUpIoYrxhYO9XQrzS8ug6ArxrM1IIkWEGhKmBdB+t57TVf0U9AteFSaXJONDpOMP0O8bBH+TTHWxtcRRV+ubm4RaTVGjX8VyqPN4p42KGTROhuwpER3OdHLNSc41wzK0pOZnNO3ZjjnS7/oRfzK51yQEFWuhDRnud0teFKGnFweMDX44ivzp/y/mzER5+OuLdzhbcPr3J3t8dO3MXoEvwCfM5abEDb7x8euvplkyW3WXUNY5XBcm5wXBUEalQrBCoULLKVYuDy0BDLgqpLGqta4LZA4CoGp/b/S92oBhrfsSDVa3iaSHwhpDMqX/nug7sCbcLvdVdiVb9HVVXQQ6MA1FZrY8K1hWlrb1b3QplQ0EcMj+clHz0d8c4XjzkuxhilOezscHfngMN+lx1v6bicxIaaAxbHTBuOdcxnDv44nfO/zmb8dVFwJIpRFLGMI6QTY24fMnzrLr07V3FpTIFQ4lZBZRvS5fuuNiKrFJnmp8cHy18UTgtm2EcP+xRGBxWpittQVUh1hd2ssrTk4ir7vmnTSv7x+esKgQLfLNkLZ12SsSFUPKSl2DqpAi7bkYQSpNjLnl3xY9QBCBEAbaHqQZUeSh8ieze0z/VPFxfItkV6AXxpH/cXz/BNAYewAS5DYet0sh9DI/6+t8J3eeYXfpZLbvJ911hobiPh4k58gPHTlGx3l9F4hsvniC9bcdGyBZajYdDBig0WmxOIMkN6bZeb0Zucd3vMvnhE8XTEaLYkVx5XlExOTjmfx8wGXd7IYg6MZ2BLUmdJbEnkHFcUJIMevSzj68mMh6en/GX8lJPZOV/2Brx5sMed3SE66mJ0irJFiA/wBSF1sN2pbhttDq60frQLEdnqY912zoN2YOKQUSCGxqduVXDBebcS4g139OGZXEmTqih14Fgt8SrYvm1ZKipEwq8eufHXV8d8qCTYtExuQ3WiYNN92kjYqtJfdV+nDQ5DaRVnk5y/nJzw0dkZXy3mzC3sZrvcGA650etyoDU7riBxJdo7HMJSG+ZaceSFP88K3hnPeG8843MfcWJippGhTGP0Tp/s/k2G928SXR1SJhG59s1zNe5euWTt/YDkqUAf8cSDAfGgD0mMUw18uoL5NwJRfQsjf3mNnm+yJ57/TU9L+G9+vTne/uYWWVRZ+Wv4sfhmW7zs9KMgAKv6+oEuQzmrTP+wcSqhu76JFF7Uqg1qrQBXzByhavu7mj8nLWHUSr1ZdwKtP8z61tiwtep7fOdjfoWM+IBsbNL3gUSsoy/Pp2enHT3jexv3bO7NRouMWjb4Fzu2QndWjTdrX3QpoOKIZH+H6OkptshxSxs6zcGlL940r6v7yFXGa6kVkkWYKwP66g6mlzL7/CGLh8fMJ3C0hLLIyadLzouSB90Obw263NYxVyiqmgGOroNICakxDLpdDoziZDHlfDrjr+djHi0XHD6dcLi7w61Bj700I9EGZcNiDSBAXVq4fuhqsV4WSHvZpNWGfF0PX2DVl6M12dqvBr4RwivYRVpWY/M4tfleQ9xbq+3VqEa971wV+6Caa1/Anf3maqp3ZOufhFx+pzROR0wsHM1yPj855dFkwvF8xqLwdE2X+/tdriQx+0nMUHs6fklqw3ULUcyM4UwbHlrhw/MJ70+W/HlR8pWPOdMx81hT9hLiwz36926R3TpEDzu4Tmjs4+tXr4VrheZs7tkmQHnjddvTtG3q2p+3FgzylTtTVKh+aRT9vR2ifje4VyT0RlTVvK7CAPzqLi2md5mV/izr/YdWdnzjBtp8BniWlb3+XOF5Q2HIVRGkcCIrweRr17BfKcBVHZJ6vDbFBw2uIJXy1wS2bmyAl4t+pBiA1hD4zYPNh/B/ocqRbZ8q1C2VfXuTNZ9XQr3mKQ3fq//QqGTtaa9bBEtzrpdQjaw+a1OAtwVT+9H95jFWwp2177arR7UXoV+/54Xlsn39tMfoG9Elp9fvcZli/CKXW41l9XljDNrXv+xYmy/V12wraw3UHylMr0O2s8NsscQWBZRVEc9LlJnVmmg9nARk3CvBKU10ZUA31qjYoJKI6cMnLM6nnMxgmeeMFiVPygnn1jLqpbwWGw51zMAHJSC1oU98Vwu73YzTLOVx2uPhfMbTxYLjJ+d8vpjxYNzlbq/HzX7MXiIonaC8QZRFXO0HrysKtlhOW5HdNhENl6/fc7PmQDXArh6kahLqqHx8ELLNQqjP86vrV4LuUmupRhKaa9bPVGP/rO7V/mq7L8HaPTXeRyARPjJ4DJO84MlozhfTGZ9Nxnw1mpFbRSfOOBh2OEw73Mw0Q3FkOIwtUD50ECiUYawVj73w6bzkw8mCD8dLPis8jyViHBvKWGMHKcmNA/r3r9O9fYgM+hQqVJjc1lBnG71InOczacNA2bxU4+LUiqjXJd0ZVl3/VGXsr5hRZV9dhL79lg/fMxrw3dGFbWrSt7zKtveX1octTL3ZVvXweIIC1mZQvvVjVQbg+x3I74l+tCDAINZakbwbaGGbpBrlRiBWg7t14T/v1h5qDTHcTtZ+ryMSQlBgtUGk/t/q+drCv63HXPos7UWw8V1HXYgzHKlHphUd0dzUU9dAeNYrXr62ti705yzFdofrF121W3nJphCvNtjamG05tr4RW+ugmYtwgpeQs+61IR0OyMcTiukMV7r1Aa9JLlpfmwzJAbkSfATRTvf/J++9mma9mlMAACAASURBVCxJsju/33GPiKtSVWaWbDUKYkFi+UIa9okP/FD8SjS+0owvfFkz2hpgS3AN2JldcDCDltOiskTqzCsi3A8fXMbNW90z4HSjjYixnqqKG+Hh4vg5/yOdhbU0ixl+3rL63StWb2G4F/rNwKrvWV3ecOMGrvfm/Hza8Z5tOVLPwvW06mm9Z2Iss65lPunYn+9xdrfk5dUlF6sbbm5veNVNeP1ojw+PFuzN5+xNOhatYSIuWAJcSenLk7pLZaxnbPTbGA6jA8EtUNclSI6TaCmoy+imQLyUf1/3IWpHeTHzdKY66kn4by9sfa/eUfVzsV0joAaaCeobBm248Yar5YaX19d8enHJFze3nPdr2m7K0/kjXiwOebaYcNwKB24d/PwS6pL3WFa25do2fO2U3y43/Ormjn+4uuOltFw0E+4mHf2kxRxOmLw45eBn7zF/8QQ5mLAxwiC+nOr3Bwj1Xfvp971XzXz+pIkz6URCAOKkYe/xMc3+PGRUVBRfwgSLQpW/Jts082Ab/v/mGvOAMqvvrgxbZmFXOYAkxhIYKAzPpwJXP9pp/IEAgJIjUKg1AjNSwrKyAnhTFQhVqTKCwoLVrs36Mzu+HJr2krIJsTkTYevwS6m0LAHEvHNv6xYZpXs1wAhuCR13UqAujpzABzHn2vAwcj0h9ndqF0lbqgetqR9bbSWG/y6SrHj+bqm++50CNMYWmtLoH++eVAeqeML4JwcLJod79Dc3+H5A3UN8OQ7wfDhArZ5zAmqF9nDGbG/K9OSAV4sFq4+/wL265PZ+gx8s9/2aN7crvlj1/Pn+nH/76JCf2ZanIhwMm2AJ8B673tBZ4aC1PD9ecH0w59XNPV9cXfLl6pp/PPuG9szyk4Nj/vTxY35+csiz6YTGehrZIC6dMZAE51AJn23hWY/NlmlMTD7HGKRNlRqKQjdPXBLs9R6pZ0zGk5wj9tP3Mmus3knm2toisS3SJPRbQjS/mnBiX8+EjQrn6w2/vrzmP335im821/Q49pspLxbP+MXRMS9mUw6NMNOBbr3BMIB4HIaNabgxHZdmwicbxy+v7vjV9S2fbjacS8NN17CeNDDraI4PmP3pBxz/5DnNoz2GiWVtgEZz1P07g/seaLq1FhAFsZTfghVybKV5eK/MnI/fMEhM+1Nca7AHC/aencC0jeWH0xTXBdmTS6eCEzqefbdzSOO4hn+O2f+PGQT4+7xbV1sMW0VjQLlsLVFFp3FPOOIx2lVbydufgjBDcazgQTOqIfulvMDumfzxXD9QHYB47GjkLypBIOezUipl22gwxeYFUgG1oDajVvFhEWuEqhQfcrixRRxiCGeZS87/z20TIMX2+US1SEj/r9VPqXtjNXYMEevgmtG1hSQD0Em0t4O15La3UGolBB6IzfTpmq7zO7/n5h19iEj0qSepLzp+fstnKNW94g+o3q/ule9sf3/cZ4nWJCHmXHcN04MD3OE9y/s1Tnsav0Uj28J/vLyjQXsBbxWvwiDQLiY8/pOP2BwecPP519x9/jV3FzesjLB2A/fOcXF5z1d3a/5yb8Gf7U34oJlyIqGwTBer6M17x8R4pkbYO9jncL7Hk6Hn7P6W1zdX/O7+lrdf3PDbbya8P5nz4dEePznaZzKdYNopRlPVvD6k36X697mEdiUwHlSIi38aCEF3u8YfhW+t2e8ASw++sc2M8+OxUE8999sWLSEIezEgLdCG43ltixPD4Byb2yWfvHnDZ9c3fL1aceYHVsOEg/kxp/sLns3nPO4mPPfCvhuY9o4Wh+rA0BiW0nBnWy6k5euN8sn1Ff9wt+Tj3vMVcD6Zct9aXGPh0SHz959z+NP3mDw7gsWEdSfhZMmYsZBnZMu2P75XD7Cm8T/gUqKC8FAAA/QCXpWNKHaxYP/xMc18jrNNPnvggYdc0zFZ5HUTdKSrJPtNUAa2hVo9rqqjW9eu/tbvyB/Mh8pcj7Ig4r2aO+wM267Gh+qOJ7bv1LStRW9K39ZU+Mpg1GCS66q+PITiXz/O63sHAF5EXdJ4s3IikQ+E08VKrex0CIiQToNRA6KCJZQOVe+xJlbyM5V7QEJb6crmrhj4l2R+ijn2GsGHV6xPdcx1vIETOhlJUTIhZCGbg0fIEkciwahojpEC/84ASE0bMPPHsbCXWCehNlMlV4WNmzTfg1j0JXQ2BL2EecwAQ2qC3r12oaBLeqD0x2g4YzyXZI5Ap8CBNFrNz9dOD0iB4TEZL1qca4BS0uK1oKOMrovwD4pmeLibzXAH+2wur/G9Q9VVsmY8yPRuLdpyD+PCqgbmCoKxlu5gxrRpsNOOdm/B7e++wb2+4PZuyWbtuHNwsfG8vVnxu2HgT+cdP5+2PGs7jnVgoUrnHY0fmHuYGmFhGo67luf2gPNJx9vVHTf3K242a/5hfc3nq3v+8eKWw/mM4705p/MZx5OWadPSxDgB8QMiA+OjiHcx3l3a97uuKtc+03daC8lzlL+3DbgfWD3HzDq0GWMBjEVTUJ9M8LSsBjhfOV6t7nlze8f59SWvl7fc9Q5oOJoc8Ohgzsl8zqNpx2Fj2RPPwvkAtoiHHJmOGyznGL7shc/WPb+9W/Lp3ZqvnfLWGm7ahnXX4hcTuifHzF48Yf7eEyaPD9F5hzPgrOYYnnp6x7t0e07SFNb8IVLedkEexpA/t5msBanVuGeNRL4Zp95MJswOD9k/OsbYNuid6dktWqgLYmUhFnmlBKSRBaT3mXkVvqShnsM4jG4HzeVhF4vD6J0/EAwFZcrvEP4OMDEeI/xmtiZXIr8p366Y9c5vQdonYZpKpH/ie4E/Kiam0Y7iAAi8w6un58d7/TB1ADSRGeAUMyh28DS90EYBlVFW+n8RnAjWGszGM90MtOsBR9DIAJB0blilNVbmbY9iGOgGh7Ee3ym9CI1XBlEYPM3GM1l7FoMiQyw5XAUcQqiLnvKdFcD7mAtaiRBRJB32LVEoqk+UF/sXqtXtMl1JVTktvZDLG+fYCRfrFUiV3VAHMWoGI4ayiQMwlVBjPfGlHPBVtLxxGGIYfY4crgo4Jc6SznioKzQmROFjap2SAMB4v7dawEkxU8b1lNRu2GySQdZYwIXjYgl16J1iga6bYmcL7q6XGDdgfF7FrRkfh5PWICA/kYeU4jSEZtIyP37EzHbsTabcTWbcfPOG9fU9fa/ce8/1MPDmruesH/h63fLzzvLRxPLcWg6tYarQOaVzAx2OOYYj0/B0NuNyMuXttOdNv+HtZsP1es3VzYrufsnezTUn0ylPJxNOpi1Hs5b9zjK1Bms7xGimhKwB+XgYTxqMxtS5VGsg0WeOvEzXdpXCd13170kDEoKqHLV/geACjOsYQbFKqJqjKjgP643jer3kZn3Hm1XPy/Wa1+sNV6s1q8HTdFP29qc86macdlOeTIRDC1PjmLieVkG8xWPY2I57Y7hS4WU/8Pm657frgU82PZ+te1474abtWLcWFhNmjw6Znhwye/8J3eMj5HCBm1hcTIe00XSc5qPgym3PcRH2DyxkQqRxfagp7pKGUVOvnQ1eCpQOipPgm5Z2vsfefJ+FafEbT0M4iV0lnMmw62s+RsKbJBwzfyrPqEistxLjuDTyKtm2KyQO5B9+Kz8/ViSo/vYuKqtkOokHPnwmwBwvEnspmKhBBJYsmZcVNSTFvyS691GRCbyuxIRp4PMVoDWUbWNVmXloNo5mUyxxYcv57z074v/r9QPFAJhidncef7/Cnd/A0iK2MOhE2mHRIzOxBnPvkdk59nbAdDb/pDkdsCxOnean0VSqbsP9fMqbvSlNK0x0w1o6zgfh/maJv13SmI62seGwDEATYlUw2IhgQ5vFKV+JEPFIEmBJQO70/7jxBonM1/hKkOe80ipVCheYaDSXpIh1NBWciEAhl2cdX4pgqv4Fue4RH+dQFBVXrBtxp6Q0PFNFQeYUmmjJ0WStUZeZh08aSh7VFkXEjLTRc7l/oUserTZtYGblShEiiuAwPrQ52fTYpUPvNgw3d+BcZFg1jSShnqwqmerKbG2heZFwqkWyGk08TPcOmJ54htuBm6VnGHoGa+gZWLkNN/c9r5Z3fNnAz+YTfr6Y8eGk5XHTcGg9CzcwcY5OHa0Lx+aG1ME5p7LP9QAXqxWX99fcbu64Xi+5vL3jS6ccThqOF1MezWccTWfMZy2zrmHSWiaNpbUNEysYF9MJ1YOLR+bG+cuAwPhQB+A7rx3aUubpQs7xj2cOQAOmLvoTKu1tvGcdjyPebDzLdc9qveLqfsX5/Ybru4GLjWNlBG0sk7bj8eKAg9mUw+mUg6ZlX5QDv6Zz63AaIoKqZS0T7qTlShpeeeWrzYZPbld8erfii8HxErg0Dcu2Zd20aGeZ7+9z9OwJe4+PMfsznMLm7o5hSeYHBVQlcB6FsshWRH0BACm112dgDH9IYRhVn1UACPswblVAMSY0ahZz9uZ7TK+WmM1bxMa0v2ovme3+IaWQGkmr9eW5BOQJVTdzzFbWhHfBZo1KTz1LUchKnI2Kd0pG2FUmV2pLK8ieU/Z8mWgprNEoIAZnAt/OgIZiXRYE62MfpZqHHOztg5taAx9ypowxqVTpSvFoImHrWAW5vIWLm1DbJimQijrv+DGbAH4IAFDiWLzBrz33r69423yBTmzW5j3bpSqDIFRrMZMJl1+f080mqLVZ+00njI202CwwPcqA6MBaHU3bctVZDqzSyMAglhtnOFsOvNo4bk3DxtgIKoiLGOIDjDcpXDELdScxvzZunIAwQ40tFR8qcgE109QqInpbATAuAgCRYF6vhF/JnihXcGUEhmt86IuXkjGQNrKv7OrGSzz9s6QvGRdHJoo3aRwlZyNpHA+1iKTl+cSRRuMN74Y7Vsez8M7nfAAAHo+P/pz0bv1ceD3MicY0M+sDw7UKpnf4m1tWV9f4wY0qRSZQFywLiqt8oVoFsRnN+SHx5/i7DyfeNT7W1OnTvFo84XS63rTcIQxiuXYbvlmGanKfrHr+/GDBn+3N+aDrOEE4UGHqodFQaW/W90xl4NA0ONOw3ptwt3fMbX/A2+WS17f3vLm75TO34f+5OodLYSETjidTnu7NOd2bcrS34GhqOe5aJtJiDVjjMeKDu0AJbpNchEcLIoN4PxFQXKsH+f3pflrPUghITQva4LVBpcFL0M6cOu6GgYt+w/mq5/zunsu7Fa+ubjlf33Gva4wYDmXOwk54b7bP6WLB0aJjr2voZMD6Aet6Qtkfh1EX2hbL2rRcSccZli83nt/eLfnt9S2fLTdcSsO1bblrQvqfkxRua2hMg1G4P79ifXnBYBVn4qmIW3EQkrWPJIiihBkJ2KDs2OhJ9xm8Kg+P7333VZSZBD4C75NoWVQjYKBb7CFnF6ymk+hKMeHIqQdaOnm9Az3b0W4MGq3H52qSaVyxIFPUlktOvt8ijQIEyhjKl1NMVzpq2sRTJFUMLoF7DfxctMpLEY9K2MdW0z1ymrWNZ2q4ioa3LRQhkDwcKO+MPqTnGPIXYF2TR7EraDHNVQIfnRq4X3L98Zf4pcvFZ1QFr6LOyUMG/iO5fojTAMHYzEB147h/fcHq+gpMMTrn2ck8N0koAbHcTVok+eGEUnWsThoHionJR414wGjPV17pFFo8hqCJ9GrpvTBg8bbLQTO5IzFAsPRHRz/nnyoLQIlfSARdiqeEZob69XJlQB3Gm4MjIsDY/m4YuhBOmYuMV8j+8KKsbPUlByTE8eTCMr70Oz0HW/cS9E19TnnidR+TFrg1ttE//Lc8F/slUSilrZN3XfWwkIV2CigSBZxHXY8fyBaNMmmUseF37MrUJ1OvWpmrON7k9TBeGDYOP6QStoHpDwShtGk6emPZ+DWr9cD5myu+uLrhJ7MJP5tNeG8y4bhpWKgyV0+njkaVxntwPVNRZsazZ+Bgb87pYo8rf8yFc1ytN9ytNqzWa27WS24u3/DZlacVw8Q0LGg4bDqO5xNOZh0HXceisUyswTQd0jRg23CioFUKz4xAMs5pLSUKP0wL4lEXfLDqNP43sOkdy/6e+43jajNwvlxzsb7j2g/c+Q1LHeiBQS3GtcwmBxzPphxMZxxPJhxgOTQNeyJMtWc6rKPgC7q4F+hNQ28b1mK5VcOFg9/d3vPpcs2nq4EvNp7XXrlopixtw8aEg3pCBHGoJKjDmtu3b1jeXIIxqPgYtxOFxHZQcKJR9Vv0uCX8MoCMOmQimMr3XxkURpptfibN/wMxHTdFTGuSpsG0FjHhfEUq/3x5p9B8uqsja0Rcc1XGVoptTrUt5GvZloJHtxQChZFpIWdDVO9m9lr4ZWEp1XNj/WH3vZ28R0LbWvFDqR6W7XmOr2/dGrMgKcvqlGHZ49d9jFWSUJlaxIuMTJc/qut7BwDpqBPBhApgoviNDwxzFzDKgqciXKlMcWmDbNNhzhOk/JA1nIGND+ataIkMGqUavEbNxdTFSdJltrr3LSAuI+Tq38DDk0G+jRbSrk8+2hSL+xB4lFfMju9u9XNXX7IWk3ZeouT03ZriddyXPPe7dlrl63vw8y7O966B8R1ztf1d4hpEM6E6cpBZBhZmC7REmnmw7wOwyu3vmr+ab43ILjHnwPidCBtjEd8xDMKtH3i9dnzR3/Ob+573ZwMfzKY8n3Q8aVoeGcvCO+be0TqPVc/UexqBqSgLYzmy8Nha1u2MzXzGauNYbTashhWrfsOyH1j2jrfOcSH3fLW+Y3IjdEZojGDEYs0M205p2hbTNLTWYKwJlXtD1h3W2BxM5VXwqjhVvNcYRKt47xncwDB43ODo+w2DW+O8x3lP75W1UzZuYHCACtY0LLqOxaRj1k2ZW8u0tcyalrkxzI1lCkx8AEMtDonxIoMIvbGsxHIrhkuEs97x1arn6/WGL283nA3KWw+XYrhrGjYShL/PpqiwprEYNH4Y8G5DXSynXMkiWNOlDfSV6VPJ6EkTH4hAvq59sot/fJsgS+3VDwuUqo4BAGBM4LOS+mtKY5n2Y+nkUfBb0rG3rHjvYnO6vbd3W/9GA/HJSrgNmOqxVW7CmvcoAaRlMFptxSQedt1LckPreQ/xJuHnwOcKNtjudyKTCgjsSjlMv+cQLYl/z65MRVRFhm8RHP+y1/cOAGwJjSsLJjpaiFF6Vxb8ScOHdNyokZS3H+4HwGhQY/Am+nDEIxr8wxYNJmS1iM0ZnIQCO4k4JdTKjkRXx0TlTIJgd0PeuTPSpdXfEiOIISixvZJJmr5RXzUhShUBD5VHbMcna2GrvDPKW2MJIkmBe4TDmOJGDmbh1A/NQTHp3zlKOF+71POQOZFOJaufrSNxx9zuAWfIZkat5HARv0mzkrIxK1O0xHGmuBKv4F2hK9HEHHwOOHwAbrwpNJbXfhsQRjuBVMGW1I+EVWskWGnWA/QD3HvPuXN8vRn4YljyZN3zomv5cDLlvYnltDEcS3BXzTB0xPLG6pl5xwTPPoKaBm8tbtrRTzrWfsH9MHA7eG6859471t6x8RsG37P0A7139L3i3RovjkEMWMEagxhBxGPFY4xijMXEsXlCfJPTqOBonkKcD5kc3jmC4dzRNdCahsZabGPojOHAtkzFMjeGvcZw0Fn2GstUlA5Pg9KqQ9wQM1vi/hRhkIaVGO7FcIty4eD1xvH1esNn656vNj2vBsfbXrlvLOuJZWiCGyVlyhgBMWOlI5N7orsRhQmJYkUrOs3nIaQWKlqPgDwFpoWHKo29fJUi0JUHJea2aL3uoYhgxGCSKTvXcihUV+5oXKsUfFz2bIlal2LxoepHSj8k8YHyfKD5LcC0A0yLT+1LFLpbZcsi6EoZXCPPStyTOUtMiyEhhyRV93y1RAUNuNxwzsAyQaCX1U6zZeJINb+TBrMTAKRLLTpAr55NkvVxGmOg9L9OAGBMoxIqI6iIIsZjRFnMO/YPZjSdsh3VGaY5Cf+4mUQwIkzbjq7rsDbkDHsRZNIxtC23OK6GJYpjbjx7VpkbmOoQ/EYKJXAvBvf5cDSpl5TuVXxMiaGnyPsQaLK9ju9e17CHFElaaCQILxUR52+8Y/5Sv1PXc8M1CidGrRb2lSJxpbxQ+qUhQCgJ1mA4ietgfJl3qCL0YyzECACkPyOyr7TjFEDpR5smgLJQZrnuU+1npWpdw+4xiZnVJZSLME8xDjJirgVvOg/rdc/9ckMIhOwoExcjdtO53sltRPAXVtMf4MSIR6bvRuYZ74hIpKX0u8HGykWb5T339/cs7+65ub7nfqPcDMrZ/Zovlhs+bda8mEx4Mml5PrE8m1hOm4YD0zDHMdGBTgesKq33SK8I8YAeY3GmYTOZsJkFq8NGDBsPazew8Y5+GFj6nvXGBxO98yydY4OPFjGP8wOOAZcAWHSTeI3ZMdGdZ2IRLYswkYamaWg6obVC11pmjWVqGyZNQ2MaOiPMrNCJMEGZqGOC0ulA6zXXN0h05xEGGwr3rKThJpr43/SON/3AN+sNL1cD39yveOUHzo3hzlhWnYGpZbo/5/Bgn+l8QQrKzRbHkbZb04vJMUTF4GjzrzWdhrZ8Xveyj02kk7KPtNKUy558EPa2dY02PCEjQEE8bWuYTlu6Llb6k1TTwcQeW1zY5RmjaHb9pUqPhnASW+QXObsgQp/4oqjG2iwm0nf4hkiIn9Gcrxv2aAEa4T8T50DEx+Bh/yALqoQxVwAgzzHFuqFbkGrrXnlOSDxL43hDDIDNffeiec1SgHqskbhdHi6uVpIdtQslghtaVivH2ctLPv/da7wLbRhQsT9e8z987xaAM+DUIxojj5SuM3zw4Sl/8d/+gtmiIVc0g7iYCY3ZahmEtmk42T/k+PARs/ketunwbQOLPe7ahk/Xd/yXqzPQDR9MDT9dtDyfNCycC/5UhHw+uYL6mNoWtWGnZYOWxU+6TyL6CopmVL9j2EnIKcE/Lw8DHN+17bfbqZ98ADci+E/BamFTBJZtYyDhtmlPR+leNYKv/L5bYyBvnMzuQHxkEpXvPykAWs1XBjuVgE6bL3JOeTDridlBDgsc5VKH7ZV7Xw8xNmWMAa/0w8DF5TVnL98yeEVoELFbTFsiMNJ6NA9WSLxk/pLrLVCBs1H/0++GxgTBcn19w9nLV/zu8y/53Sdf099uWPXCxgk3Tnk1DPy2X7N/d8/TxvDhYspP9ue8mHacNoZDY1h4WDjDVB0tgc1ZVcQNGHVYEWaRSTuThFc8RKvrcNKhswCeB5QNoUzJgDDogFOH96GEqUdxPgD0UEtDg1vAGowJ4NmqYMXSiQ3BhhJS0ESVkJAXGazvaZzD+JCuGfJqAlS0MdXNidALDGJY2ZaltdzScKGWl4Pwxd2Sz2/v+Ga55KwfuDWWpVjW7YShEbQzNI1lvj/l/Z++4Ke/+Ignz5+F9TEl4mOcEeIyDRuaSEs+ewMsNloWS8ZPiQ6pebvJ/5KtPxOJKnW4sq9oJD6vZUdq5jU+shkFeowRjo72efRon729eRBZOlA4l9CIwYXNHtOBS4c0H7MMkgBABEEP05PDu0aTdl02WuCAtXZS8cS8eyRWXSUof2Y891vpE/H6rpMwx9fuJyUqXoRexlMmDU1hb2kPxz64EHocJU8te7a+p0P4qiR3okG05fx8yX/46//Mq7f/ntW9C9UBY3kgY+wfNqgf8Pr+CwEZ7xQGQbQRmE1befHiMf/2v/szFvsWJRBvFiY+Gm+Tv4ZAfBbD3mzBe0+e8/6L99nbP2JlWm4by+/6FTeXbzi+3sPqmg8Wln+zP+Un04a9wdFmAABZFGlC6OG+p06fi8QsdRx4ErRV0Ny7AEC8NAOAiPhzY2OB921XSrvJ85n7V4aU6geEzAjF48txK9vCSdP/1WNJQn0HE9A4jhQDEJmA5kDHsR4TtKjIdPJuC3OQ51Zy04UzbqVHpcCp3MO6DkDaePF/PiL8NMdBKw8fGQbPxfk1X391xvX1PT7WUUhdDDGbVakUCfQmXvMYFGJUss1zkLr9DvwX84hjXzCIGob+mI9++oy/+G9+wZuvz/nd59/w9VevePP6ktvrFcvecuvg2g9cuoGzmzv+6faWJ8byZGp5PLGcTAxPZhOOmxl71jBHmSg0KJ1zOWvC4Om8ghMk5otkQBfzpb0o3iiDEVQMA6FwSZhHAaP4piXliGcdSaLlQQMo6qxinEMGj4mpZJoCRhNkFMXGFETFoGLpxUahH+pzrA3cieHOGa56z+vrJW9Wa842nq82yhsHl8ANwm3b4NqO3oBMDLP9GcenR3z4/jM++Og5py9OOXp0wGw2AXFjAB6Bs89QTUFjqmuhzEBdIjGf20Sa8RgaFIfsoIBgWg5EM95KtQsyRpxHpSibpivAH8+zJKWrCtAY5eBgwdNnJzx6dEjXtYDbilQXjBG896Pvlm4WK1eOdo9afD7z3pN5n1AAgI/1POqwiFS3wxNcVEiIF9FI91ZzLD/FarL7GlXqrJSRxDceSNCkcKTOxIdlBADI3xQ1D55NSx7CU5LFI/EyGS1v6J6r+FrgQ4YJb9/c8/mX39C2ht4MMWdYVcBZa3609YC/VwBgrVXx3hk1gzFh84gobSvM5y17e23sQpIICYlGJBwlhEpg8E2rdHPD3uGM40eH3JuWHtjcDdzew2be0aG0+x3zgyl7Xctev2GiPhNq+kbZ4iZuiYr4opAqfqi4FbLwDhpO1mS3XQNaiFXiBsjVAvGBOL/N9r91jdnSwyudXpgAgEaG/53talO1GgWWGX8lmcdMHgdRAPpKqNcb8eG4BFuEwSgIqTwhardeKimX8ZH8FfHRIkEwyzsxWF+h+sS4Ae+U1uxj1fOVf8m6j5ptNAMGN00dSxC/8uCYN8lpXaUw067hJrNvAQkm0k/XNcxmloP9KSfHB7x47wmvX1/y8uwtX3/zilffvOHuesmwXHGzEpaD8NY5XjplbzmwWG/Ya+D4bsOTdspp03DStJw0LYfGsm9gwU0lGQAAIABJREFUJsoEF9PklBaNtcpjdTQFSwRW6vHeRyZQNFxNAFETECOrpqlCetF+Besj00z7I74frAiBJp0I3rQMKAOWtWlYYVgJXKvn2nnONwNvNz2vV46L3nHVb7geBq483Kjl1hg2VnCN4FqY7nUcH+1x+uyEJy+e8OTJMU+fnnB0tMdk3tE0FmODThdJKq+vQXMhnEJeD3dNGHYpQx4aCdH2ISYmPVeqUiRK3TYkJ3e9YosyIh7URWtZmmjJgNZE15k1wmI+5dmzU46PD5nNO6wp3xtxh6220q30XOF+iVYT2JC8zjntV3NIcgQt8Zu1CT2O22jQsIMwTfsz7dWQgpf3TepLDJ7OYQxaPpxv5cDmaozbwYLVghVFrebpEQCMvgHJqeniN4xqBgpSN5p71JSmfaAtoeH+zjJphQYNpeoRrBhvje2ttf86AYAxRrXXXtGVFauDOlEdQqTwZgVqo+8pwOW8GSMyjpwYcIFBywDGIUYxBtQKK++5cgMXw4aVSVmDgo0BTUZCrmkpshM1mbxBfDTjJsPzGH0WNVBK8kFE94VhhjZHiWNZEPn4S1XIJhfDqIlaEu6gEGz8V/xowqWjdyv+7CWMfxycV4+j6lx+rjxjspZdMmKT28PEZ0OKq8bNnAeaxcfok/l7rv5HGV+lIom40Eoyk6SIfmLOcsXngkYU/xfnxpgCgpIwF8BaYTZrOHl0wOrunreXN6x7hxcfxpD4+oPCDDucAFkLjjSZvi9k14po0q5q33DU8oxHDDRWaLuOxd6E48cHPP/whPffnvLq5QWXr685f3PF+fk1N1d33N7fc79yvPEO43ua3rEYeo7E88hYjo3lSRMyCI6s5cAaFo1nYWFmLDNrmKjQoTQk0yTR/J687WFMAdtVaxJyd8I4lGI1qf5DQmVOERsTbE1sKaSiDXhW+CD4BVZeuVe4HTwXfc+td1wMjjfO8cYPnPee87Vwp8oKx8YImy4E82lr6RYT9vanHD6a8+zpEcePT3j87JTjJ49Y7M1YTKeYcDJLUBwyIKn3VhHVEtcoC6BEB7U8rSlBktAuNTcCu0qCNu2ch3BdorYvKQBNQhErlaRVpgh+iVap4J6wRpnPOh4/PuL40YLp1GDE5X6FMfhKyUgdlqL1Vq7ossK++nfav4m3yKj9kgOkuQ5LUqpSfI6JdkfLFi+NYjZ3LwEhqWMjgqu0zmKS2J8UW1DzStkx1nrRJAv5upKiRlae+FyIZQlO3qLQZDd0bCPt5YhVyjdTO+oZ3Ia+X4egI1VEDGJkaKxs2nZSn+L1o7q+VwDw5ZeNPnu2XinmzhpRN4i43nF/u+T65o6jk1leFCHkIXuI3CYwJUVHTN5ag21MME8CK1Vu3cCdHwIjMiHiuJHgWwxtBOESrmS6T+lzVVR+9DXnPOB4SaUZ2EwOoU85FFpC7a209X1CCnnbVKBGEouIm0PhQcSwpp6F+aj91QUopDsRvVLrplI/zni/hPZV6nlJLyqj9Ka89SODG/UlPFNcG8VcKSnTIj1Tdb/8UUrXprQ9qZ4O7rntjQ7BpJ1iDMzI2CdK1OzJCl3TGBaLjqdPT1i7nuH6lt45Uq63UVf1Na136cN4LmJqaQogzGM3+b2kWQVlo9r3klyBgohFxDDZt5zs7XN4OufDj15wf73k9asLvjk75+Wrcy7eXHB7ecfq/p7V8p671YarwXHuHNNNOFPgwK9Czrw1HDQN+63hoDUcNB37pmPeCAsjTE1DJ8E42lnoRMORxSitBKuR0RTsGU/gjPPi0ZgtEwIGnfgoCAy9GjwNvVo2SCiGppZBPSs/sNSBtfcsvePOea4Hx2Xf83a14WYYuPWea+BW4F5gRctgFW0bzLShm8+YzeYsDuYcnx7x+PERz54f8/6zR8wOFnTTjqYL8T2BeW8H3dX043OtjLTbwhXWVmoCzaSnaCppjEa3XHEBhjLbmsEEouN1T3SkRIReqlDWYKT0RhLxY4wyn3ccPzrg6dNjppMmAvUKBDNONizGLNmWi999xf2mmVcVME1qv7ojWv06/iNeLj+X9rxPDyULYmTA4zkpVRRAYuKFloer/pDGGW8UmSLV+mpUXKCuXaAk+4eml0tf0lykJvICx75EC6LScHd7z/XlDc5pES/qNiosF4tmzR+2Cj/Y9T3HAHzm+/7ZLbY9t9KpOhg2ytXFHa++ueD5e8d0rcTjGbUQH5rFoRLSjoJf12BtizHBbeAQlih33rF2AxilM8LUGiaiWO+iBl7azWJJPalalJLWVSr60tHmkUyQ5J5JfTdGv9Y4tVzbCTNatVJaT4ay1JUckQyjrz+4KiFVAnbCW8V6YEgFcxIYKFH+pXPBUGcfBLaVx6SK3dkeaWFuwYVsMiMLpuB6/HFEGs1u8X5aoZSpl8ufSgUjZKQLPJjPfKpzbBHxNK3l6GTBsj9i49Zsbjf5bKEEx0aX1n8qpfyxZ7wUEaTqCEJsrVfNnhO4TNaVIJDaDrrWsLd3wOnTfX76J8+5vL7n/O0VZ1+/4dWrN7w+e8PF+QW3d/es157NYLhzwttBMYPHek+36pmu0kFDG+a+Yb+17HcmFAFqDFOj7LUNC2OYiTAVYWZDkaxWoY2BixIJsUDYwKIHURxKrzB4Ye0taxWWKtw55c6FUsjrwbEaBlZu4G5w3LtgDbhTx60LaYobFdS2+NbgrAWraKxDMN+fcnB8wOnTY06fPuHJ88ecPDnm6HDOfD6hMQqxlqNKSj+N1oyd9JloqAYHRa2THHBXr33S1uubtchNLdXrraPfR9YlrXdSoZbxnfgvUabTluOTA56cnrA37Qo9JVkliapMFp9pT4z4za4gCC2UKlpZrGKjqZJGNVP5G6Ohbj2zDb5KmG8ItNtCKfGleu7TfBqyz72K7B91oIq5II5jBAhGVw3KZHRPKOPOzz1w7aZyxnF21aNYhsFz9vItL796jXM+4hRlcP1qs1nfzGaz1VavfzTX9x0E6G/7+8uZmX1jrG7EyGRw2DfnN3zy6Vd88JPnnDyeQxtzs6P/OUTmRq6fAlZ8CMJK6UeqghNlrY6VH/CuxwCztmXetrQC6BAJJMfZ4jVqCVF7rIPPim8z+oW19kGH57d9bul5I8VHrlRgtbq26YnqESUEymmda17zjR33qmmmxuaB95kIQ6s9Vm/6DBIC0k177EFSZkLUaWtKGfkuik52GxMTYTITSWbYOgI7fsOT0oCqAL0U1BfXomZgqTyxqIlWl4e98LmmQfySCRamRyd73G+W9N5zs1zFnPZIIyOUtsUws8vIUJ9hLdFqEQBW6kuyBKV5swSXQWk3L6ckdFNAgjGG2bylnR7y6NE+H3zwHje3K87fnvPq1WvOXr3m8u0l11dL1nc9m+XAejWgDu68YgdH42CigvHQrQYma0cbc/xbYGENe8YwI5xBMBFHi6cTaMXQGouJqV8aGZ6Lq+FEceoZVOm9sPaGpRfuFe4UVh7WeAY8TqFXoQe8sQy2oTeWdUOs3Q5YpZt0TBYd09mE48M5B0f7UfAfc/rkmL2DRUgBbiT8Z4NJ12d32hbtQ7bOlD3mY6BXeb4IKQi+fZ/BXBKsGQhlIRPWfUQf8Qs51E+EspsiPaS6HhS9M3WwmMdDW8bAZDbl8ckBj08OWMynFd2YLD/TfvNpnYTK4Vlo2MTnar06nRUQcc7WG+FKOVDp7w9CY0bjf2jnzrY0icGB2ToW10gLT9oqAkDeO9uMJgH3uEiJH+Xy3ZFJ5f2WmVbFu7OLOcqYFDex/Vx2iaYeJZ5o8Co4Z3j58oL/+g8f8/GnX9HHeiNt2+pm01/dXF++cc79a7UA4FvvLxez6RfSNm/WQ/9ss/Hm6upOPv3kKx4d7/Pnf/FTTk4OmEwbjEl+GkHFRkEVI9pFEG2CmdULm0HpjWPT97i+xwyOiRr2TctCOjp1MEgsziTZVKVUVSljjm/RccgCKNBA2uQ5q7OKyk9bJ5Qcqu+mzbRtKi9bTB7e0zBGT4ViRw1oBBUpqKbWKscgJmzS5FODEvgYI+c1YmshoucUh5FaSX0s5vw0dpXQfjbjFRYSvq82bqkQVe0MeB+1x1FsRWINYV7DmtSCk3jYERVDGF+S30sajua5r2zzgOIYAEPTNjx69AinDe78kuVyE4rYeC17X4swT8wlWE7SvFQCJwqf2hRqvI3j9dUSpufrIKxa84jlW/MUKY0xNJOOSWuYTiccHsx49vyE2/sPub264/Zmyd3NiuvLW85fXXBzc8vqbs3ybsVmuaF3MKxBnMmpd5YWg6d10DroCP9ZYkqfhhM0jThEEv1HC07MRU9xFj4C6kGD0FkhrCWcfRIO5I3F0WIKnoigRrCdoV10LOZB4M/nHY+ODzg+PebwcMHR/ozF3pz53ozJfMJk2tK0TVxXB+rDuUZxT6Q+ZYpN1hiRKk1Wcr8T2eal0bKOyQKV4EEAAJKzOoBg7t9Jk7K1hwp7jV7Nik8kZB7sfunUPxHFtobF3oyTk0NOj/aZzSaIMfSRxlJPA0+IQFkkZiAk8FxoLliqDV5c+X68l8/UqN/QwlPCgVzh11CZfEuOVVk1cSrJK1EJ53qOMtCIv4umQGahuGbry+e3JO/LKgkz9isFZpa1SuAw9XXMl8sa1+5KRr5+jWuah+3jmD1sNo7Xry/5m7/+r/zt//VrvvrmnMEpTWM4PXnk2sacvXr95ku3udvwI72+fwvA7cHd6TP93Bj9VddyMPR6sNkMnJ1dyN//3a+5ubvno4+ec3xyyHzW0VqDbYRpN2XSthgbNWuFtSpXV0tevjzHTNdciPBqfc/N5SuGy2togoVgvXZc4Rj8EkMoMJKYdzA0pMUujoYxCEh+7jrQLTACfDLWpySidwO7hxHidZb5rnsRAKW0nC2BGP5IYEOjDz/9UAlhNGykbFWIv1eplWMiLwzlYf9SakzyzzMqorE9juQYqb9RwPaub0TYpQ/H+12JEgnMFCtB9Y3Mi8fjB2FwBu8aDFO886zvN6zWfch5T8JYTRV4pNHPW4ARMcBsXFchXOlwEk2ZBqPZTC6AZCUpfS5ulQRFDUgTmWyEcNKwP99j3s45OnRs1gP3NytuT2+4vb7m7m7F9e091zf33N6s+OabS/pNml+NJ7tp9lnnfHwV8KGK3zijPTHIcaZMirQOwbkGLwYnEfBFwabVaNKcTScTDk4OOX1yyP7BlL39CYv5hIP9BfsHe8zmE6atYJsG9WRAgzWoT4VnootJkp82anl53xYtf6SRhy6HADINlpwc9ChJ6GkZOoKkiP0YmBxcv1VAbibGOupctv6M448CXKt+Qko/VGCg6YT5YoLZa1FvuF8O9OtYClnDOMOIitUvtGeyIcRLLPtbfd9otABI6UP4rh93N86HKaHu2X+/S/tPaY9jwZqsqAXwiIJJIGsLRAgx6yCfIrk1bxkAhDgbQUqcT+53sOymg5JqcJAfyMtTrfFIUahfGtOTEspf+wFWy4Hb2xXnry/5z7/8Df/33/6aX//mS65vVqhHm0nD02enN7NWPv7is99++utf/+pHex7gD3AY0Nfr1a3/fLJ39O/nk+nPh4HZsHbd/XKjn31+JheXt3z11WtOT45YLKZMu5aubdibz5lNptg2+ZENjbF8Mj1jMvsn1DZcG+HLzYqvlndcrJdo2yCHewyN4XPtmfoNISVuvGFTgZpSparaSCOBUTGXCknaynxVvxEYDYwIqgoayYlWMhZ+5Y3Uv6QJ1lpo+NNkjUFzVoGM+kC8VyHlbDIv+sODPaZpo8mof2VkpfBONdrSQDKLS1WgJw89PZ/mFIrZtvTbVH1O3XonBpCkyWh8N4KB7SjiEbAJYhcszgurwbNarbm9WXN/v6TvY0GVeEa91zguiQDAVZEp6Xx7X7lskljMYPPhuiiACYLM0MSMlwiefNJck1YmiDSU4EgoJ0raULpXhXAglGDslOmswdsJ0i3Q5hZ9c4NzKUeSmN1AVLnS3kqpqSFo1tRBUhqKCGUSAZCUtlbFhkt0OUW3U4jGrBhtAtTtlHa6oJssMI3FOWF571ivrnnz+grEob7MeV5jY0I+frWmGaZmoaHZepcCa3NuuwhiTOhiTOXDuy0AEEJ8w5ZPHMOiJkb8p325LS8QoIEUVLuVTpitBdFdkU8GjHyoROoPTGbC/v6Uo6M9uomltUITv+sjkEmwLBGWF0XVBAuqMYixePElM2W8U/O+CvciD8kbLSki498z3Y+e9TkjAKphb6VHAlhNHCQ3M+IiBjDGRqtTJZRHtUaCUjPmCUpy2Jh4fHLofNn945HHv5cHq6YSv4/1PjI/CW86r6zXPefnt7x9fcnZN2/51a9+w9nra5YrByraTRo9OTkYDvZmn8ymzS+XMnzGtmf1R3S9k7/+ka/pez/5kz8/OXn6P5+9vfsfb26HJ5tBrXMq4BGrGImo3hi6pmHStjRNRO7WYmOuqHeewTt6A70VloSjLzEC1mDiYSozP2C1z5tNowaUBE9GnXEfPRDckN/zUvLEhXTETNlSwT8aL5FROybluKJVHeuSc50adRWaTQyjPqEVCVSUjupNojM9G6qwR2EoUp298YBbhbYqQJPPUVIffIV582goiR/3S9p6Ln7XjL4R51hieWXKkcMaojijppmeK286CcDJRoASgFU4Unl8lHD8fgoMTLOvhBpf+o7xbg+eoJ94DNZaem/ZbHqGwVWvJ8tTErggLjKnaKUMBWLSoga3gVGN4nocZDn2jWoQFmop9Z5DSlhyMZV3DaWwUdGeJL4brCBjpmisxViLc8rV9TIKblMEfp6m2ru7fXBN+vuuQ7KSdinkym1aA4AIDEYAIIxKRLBGQQZUh6pgjc+/Z4BVgycfTsgcZedEupJox0jzk9NGpSynMRKtBjGiPHrFS9qjZgkWhGwCBhCqXgZQErDNGJgHYrA7AcC2q8AYCdwijSO9iyBmwDZK2ylGHMZAY8GKxsj/3Gpeu0DyYZ0MghjBmAYvsRhwZCr5WG0ptDjaWxk4p/Lo0R25vfQ5hY4IBDMqjNaucR6SaNnbJvYl1fxICaiJtxhjw8mUW9+poAc5TFpLRk02wmnMqJJwVkK9/pm+6nWLCsvDAMkUZ1bRnwi9g+VyzeXlNfd3a5QGN4QqsiLCdDLxj47m7i//zS/Ol7cX/8vbl7/7X3/5y1/+PbDmR3r9ABYAANY352dfzJr2f39y8uRgb+H+h7eX98f3y970DtSpOAnL6wDfK5vVilSaViSWftUY+BO1WmcMrl48AS+GpXo28axpH0vW7jLdGWo0v1twZPZc7YQaN9ZEoqMHwr9s9J2P268JTsupv1vt1JkQeXtqyhMoqU7VlgytS0rhejgujX1OQj5rOlofDloBgMgwRu57kmiQnd+oxUhuTcLamWxWLwws9SWY8KpKBEYz8Kv7NZqv+PddIVl1X+vVq1mUGItXi/OOUjwtCqv0frSOmFTgJsM3HXcEE9PowqoFIR5naFcEaICuJDdNoM9ULa/AvLQH8mDiOyNWluR6CjSLGk4AMNHXm7T/rHGmNNBIQVWQWjEhD1RBMfGqtcIkDFK4WArykmyhKtqWoh5cBFUBwOYRhPiRWltOV9LMEqIUiRYMKe9mbm9j1lC0vkR6K7MqMRUvpacVwjb4LDBzBYQYx5EsAIoPwAPK9yXNc1qgNIZ4DHq22lTX6IhujQW4HGIcxsQICqMZfKSyyamnGl0sqWJgStnM4EUohY40leStauBX9wqYjv+MCkLyeJkMrPKCxPEMeW8HHql5XYn83PgQ32A0ZXYFM37gQ2PbbAqIlUr4Z/deIZOYYqyje7lbkTxqBaM8lvZtcZ+Usx7KU6ImP61SFCLvwQ2OYfAMzuJ9AHvGqnbThsePj/qfffjssjXub242q//z7OzsU0JIzI/2+qEAgF5fX19PJtf/cXHw6NHzJ8c8fnL6V1++fHt0fnFtNmunKBKCAPMrpFKZRF+fxI0ZCC34xVIMtoRXYoBOeMdTFhICgWqRm1lrHwuMSlgnfpgQRD0gStZqfrjqR7q2Mu0p8KEI8SQTt0VEykquDfE+s4EUjb4laCldrYHJA5ASmVfyO6dnEnbR+IivOrXdv13tP/ieFCVXqy8lg2CKXoZtO5mCS+Y98lv1+Bi9OwZoqQdZ0FeLUORGERyCwZp4r6qGWNZTML4EC6WEsxBMVWbCIDloKmhcNZxLn009jFAnT3ryXW/NAyASciXyHFRCNT1mgHTKWXJPNY0EGpM4S6MI6Tr0KdKT6ui79Yzm28llloCSJsp3WdSWo1erNiphm2IEJFp/vE/jlAoExLe0ij8QggAXCafyojlINa1jEEBa0YkUOsh9MuWXBABGpvsSm6NoNMflHj+YG83vRmGviUIIIAK/NR/VhOa4lTAO9aF0GT4VQAvrbLQW1iEAUOO8hUDpxFUijUbiVZQhWy2EpF0PtaWCGjBFXGIksd/yXFqaFDMxGk9Nm+EvxhX+KxEUWDUBxOd2tplMARvBWujHz+y4NM9NdGHEuay6VZGE5NikB+1GZhxKQEt0fyWgFPeVghiDkRCrcnS4pz/56Pnw9PGj1w2bX736+pv/4+VXX/zj2dnZ7Xd2/F/4+qEAAIB7/frLs6PT/V9++NHz9w9Pn/3s6fvP9z//4hu5u1mJc14D9VcoLVNfRLbxdMDAj308da1oJyFIr/LXRWY3IlLVWnneulJbhSiTWXtbhAYCCf/W/JmYWLOLsEbfKLp9CeTb3ZctZwHj4Dn/4I30YPoCjDOWR3MV/11rL5klVCDgXdfD2So/7AIA5SqhgumnvCFHaP7hc7sulWhlqcyqId2L8drXna4FqJOcQhXM+370eOqL8cE3GEU/Sqq5rnmiAg3mN6vvF8243EsgN5i2VesMle1up5kwmd62LxPHG0BVYmSmREVLEoGjDZH7JyMAML7y3eTHjkwU9SEmJk1UBhfFbZFBQ0Q6YyVfIr4urqHifw8PeU1ndcaa/iYBuqiZFmkSdmAUuNHsRwIAqdXRHNQuBd2mNiGLRuPy/AU6qOZmtFGUFIKm2TXjx1NeReCqgHhTGVk0f0d1QGUg19BXJMyNKcA1mE6z8I92tvy3GuqNV3bX5vBl/SIYLvgorWqeltJ6nLK6JHm+5xJA0tzPVH1PTeE7aZ6zNkQS5rFfFQVudXoUVJhpTuJB9GkAGtZXVVUrhiQ+0XHdbNqjoQR0ETNKLuYlQmNb5vM5L54/1p9++Hw9nZiLLz/+zTfn52dXm81mevrRR4d2tZKzs7MlDzMkfxTXDwkAZPHkyXy+vz+bzCfy+OnJ+hdPnrun77+w97dLhn4Q7+JJZAkVV/SZD4ysBEM5drUg3pEPkCKgwt/jc5o2e2irFo7bvv2w1iUdakx/caub+KVI+Ua3n9u+CgDwuQzog+mq/tsiznxtIWMtGQ7vFM7p1wLlq6f+OGA1CCgtn4rz/c7n0XReUBFH35UCMHpXIhONm1qDPzJZiZPe7pPlu7wc+uljS2kJ42/h8oWZ5ej+JPSpQGh8lvQhycLSmFrTosw9ZGtDtoyMxv2AcoFC29tXYsBBGoQg0aIRlxZNXJOxrK+E+HgC8r+Cth3XN6NezWckJMaYxyrB9KBxblNwZMYvKhBT0XKaXAVMw8c8qk5DPnjwnWehk6VQ9SeQj7yNfCQHte7I2MjTmlmOPPgpTW4oJR8sQQ8bqNaUrcndcqTnEsWRTxkfvRtV8G0wTafInnR0UzL8RAEfabLyhMSuJuDCqB+J/lXfvblKX0qbAhmgV/r8iFIEMD65DXR0b9c1Ol2w5hcaxmvE6G6esQsIRE6ewLgEAIAWECQFNWuWL4SBJQvrdhh1ONgsAFP1EsMFwmmAxhq6rmN/scfjx8d+MZ/o8u662z89efbnf/mX/07hAx2Gr5ZXV5/83d/93cdnZ2dv+REGA/6QAGD64uTkz168ePI/HZ4e/bvF0eLJ4mAif3L0EzUYUV/MK8kkVvPiOsgnQuEK+RVC8fngn0C52xpVOfFKYt18sh9/rB1VsCD63UsOdykf6UZCo+TZ7xSoFVImujJ2pYrlqz7wYtRI1X593LT+PoJTGKf5VS//gSCgxBmEtx7yxRBD8N0AIAjCkanx9wYA8V1vMuMhMkUT+xAe1JFpP7+vmpmUZlN5YIRB2PpsETDxEKKkkQW6iTEZtd/Sl3XLftkkBLbIKxmpQpEaX76BL2uruwLx2NHn+hsRXGJyoFZaIxvBSY2xvdS0VsZSvgNOC6jKBV0kzV/Zl+P5jb5q8dhUqqUCEMHsruo0wW0oqX0ejccyiprgryebqtXEVM0c7BYDIPIZ8ASGonmjF9pPlF5WKQgJMaaCSwVnGAEjCdrmBuMcGLxvqqEnSaMja4ak/xOHYkVMTMlEooujpIV6NUIZR2k09StKZckxQWPBPuaPaY15FxnlbqdAPZ/jrypAp5AOQat5U7IwpXffdW/nJyv6Dfw/aNgpjin8kMz6Rkf7IvcqrKl3A4hqySsIrqXo5tExaabgcElDJ8U8BWquAJ1HNDKyFKMjAtYYjLFiQAbnJyr77//kT/7sSd+v/nt1bnV/c/32/NWrv/3g4uJ/6/v+P5yfn9/whzDYH+D6oQCA/PSnP91/9t6zv/rgFz/7q8dPn/18Np8u0AGDxVij6RwAjTbSdNhr2ahCHbG7LfpT1HRCv5CAdyGH0fpXaH+M+xKzlPG9DL9TmwWWpPjSshXDVcdmh30QGUZQocL97OMjeifShpAc8V/uUd1L/TGllK5WTC2NfQc3q2evPka3jG0LZIxmpp6r8eTZfDOuUA4w3DXPGQ/FuZGaIxcBOf7n7nvJ3xeZXjI3jvta5rkWvkAOdIi4LPyWQAEmB8+JT3NVBbsVRQKIQWzJJJ2oKAt/Gfk8y7woqW5DuRcj6r9l/vIXtickft5KOf+8julPe2EEAOoJi2NJl8YYVNdDAAAbY0lEQVQpMlFYbc9ttbciu880pinGQ1XwgRunVsK7quC9mhCYqj45ar3TBLHCcByqXkMqoKpXr6qi3sdDalVCUoYPoCG4VLymMyaU8M9gBBYGEVXvg9QUEZEYwIlK8p0nCWhCCoHkMv5ixAQMICYGMagaMRZMjmSL8FND5kEhQI+KiErKzVAJR8qWR7wYURniXD6UFzVfC6QjgE/1igq9SK2cBF7lQiETDfxlq83oPc0Bq7HH2wkIorWSU77x3fck8t3SYBH+iYCsEt13RhIxRNAW8VzNw4x6TdG7amvIE+kqj6W2L47hX+hU4qZxblVRK3hBjBVtNO3k5FYQ1EQQN6i0xthmNjN+2nWwUCsopycnx0ePJqq+76z9x7/+679e8iMLCvzBggAvLy9XB+dXX1y/ufinSdO16vzjoR/220k/bdtJ1zStNdZYp95INJ0mzSkj6WpTbV+1kMuhWrIl7FJnIsYven8RR5Uo2Gq9hgThXtBEEimNC19AtQlS/2qfWpJ3tcCk/EaOuk2BSxrprn5O8nPpvbqPJe2xnqARts2dHJ2uNdrwW9ye8WPv+jULiuqhUd8qYTUGKOWzuwQe77pXPT9iYCOQp9lbM6KHmPY76nN2F2zfqwPJcsPVulEteNXRyK2l7nn+Y1v4vuvet89BZqZAnbYqses1aN5uazyX418znWZeOjZZ5fZChbw8IylJMghor6WEsuAlcNxYa0HTE4NzGgMr1XunGri+D6UaVdX7AAxUVVS9cz7c8y48OQQp7/DqQfEuggOvKWzHq6rzBBCBqiASYozAyNg+LsaY+GveYmKMCCLWBnSAWGNEjFgjYkIiLMZKCFUQCal/oSkillARMcGjL4qJSR4BOGQJTQ5BFERiIZ0gLE1aYY02++RCrwjBS+KGlcoUMM2ITkM70V4uNTfMQH5EjCrRjbRNOw9J9uG9LWunRNmf6CugnmAOjGJa6xglwUe8F04v0IQKJOLDBAfDPGlWBjzkiMk4eCMZ+EZDnUioN0FURJWYUoJG+Bdvl0BQHynKiIqC9aqIamMb11q7WVp7e3t9fX65Xv8oTwT8wVwAFxcXy2ax+E/HXx7fusH9/c3l9Xum7V5MZ/Pn88Xe6XxvfjiZThemtdPGNo211ngxMf9PornMS1icOqhnfEn1X2Jduxhe4YZ1tHD9Q3mpoOhvQR5bbWwFoO5+J/09M9aqmer++Nmtkb9DAift7l1uz9znSliWe+/oK2Ps/G5o8O73UyO1sBo9qw8e/dYP5Smpn9/1TsVghC0Z9x1jfue9d32nGohW+GFXGzvJZ0fTu37fdaX12fWLvPNfD/r3cBpr3Ur1AQioflOI5uYgtEOf0g8V204c2vvAuQfv1XuvIN45Va9O1Tuv3ntxTtV777z3AQQQ/u2c96ouvODVD94LeBdCB8M3nHr1g6pI+HD4jteqW1Huh3+LpORJgtA2ghYLcsQExlhr4mWttVastTb+JuGmGDBiDMmSEN80Yq2JGMCoMRFnGIk2hWxD8BF7CAgmhDgi8XDuLV/+lvslRMHIWOwKEkwgUmzi2SKUQWMBuarpXMCHfHFEKKX9nXcjMtlFMSPQGCyqIYTTAOp9wAIRKYScE496n3BiQIheVb0PVqb4Ib/tAymBJnF8kuZNgIDrvC/xxCldUQQf81TSZ73XZAcJ9Ck4VAfd9Jt+s77t+80b8f7r25ub/3Lx+u3fbK6uLvkRAoDfi4f/kb/XAYvJZHL6+PHjFy8++ODDFx+8996j09PHi4Ojk8m0e9Q27b5t7J4YuzCNnTZNM22btrO2bcVaixEbMbcJUc7RBhyBQTGnBQUZCuoNQjFaFSK4LTp1AogJf0fDUBW2/IApayk7mY+oZbsZEswuf63VOi38VYVcZqVsp7HY3RZ6po5a31adq0992zXeK+WFmqdo9R/scKv8vleC9umf3yV8v+UKHuSqrVE8x3a7Jbt+dy33f941Erp/wNzXIGqX4K4jNd4t2B/2ZbuNoACN/KY8UMVyA5FGZVQiJwnxoJ2qoiJ5M+R6GtGkDimuUjWeH6BJ2pLsAVGjFx+M+F7VD8Ogqqpe8eqcRmHvvfNevPfqnB+8izDAexd+dgEFeBf+8AEM5I9FM4FzHhF1qkpstoiQiH8E9c4FeeI9IqIm6Q/GZG0ziPAg9cVa2zSNtU1jrTGNWGsl/GgaY42JiCB4GYwkyBB0HGvFWoMYY60NfgWR4GJQLwET5KPLaCI2IPxAMhqUpVNJVoLwTEajolm6l4BSqZ6IPcz7Jtb9l0KliS4CU7MVv0qxB5KhwwNaG5HmmPI0WoMku+58AGnhGCAXjjBKoEzVB88OmikKF2ghUJEv617Rc+xseK10QAjeGEkuSxnZD2JoiY9E5LV3fd8Pw7Ac3LBSp0tBlkZkKcLKGO5Z97dX19dvvvj8i88/+/g3n3788cefrVarl8Dy4Wb7l79+aACw62qAKTCfTCaHxpiTR48ePT48PX366Pjo6eHx8emj4+PHh/uHR9PF3mI6nc1t107b1k6atu2sSOuNsWq0ETGNMcYIWDE2/DXA62BCQ8PmCfmvIewp+lmDe1cl+aw0bpvko0/C/gFTTtyDAjxyqk4mvgRwCzHKlmRNwVKlL2lxqnezmlaHK2r98D9bsG2D5Z39/CNdmgFAAUE+M5jveruOlNYIAEolRtGq5Gh8Lrf7PVG78s+D9tthd7WQ/3/bu9fexpFjDcB16SYpe2ayCPIp///XHSB7mRnLIrsu50M3KVrjmU2QIGf34H0AwzddLFliV1dVN5neDwDynZ/R6TqPD/EIADjuZ0hMJf5OAHDMiM/3f3QRJlHwflKg/ZydfUOoGNX+cVFPzXSjfr6+MR5Hz9Na9sE9MlPH58jMdI/wSEsK9z6uU6aHR6qHe1q0iAi3CPeeHzDzcDc3MzPrtxARnEP0QcHdPTN9ZBwig9PTc9x9EnEKBY0AIcI9swcAx7urT50pmZlFVbSUoqWUwjyiAC2sWvbMAIuKFO2VYuY+6xfRokVqLaX066uyalEVUuUU5kzmQsIqxKl9yCdmVslRVtCjgPA46z8GeOmdB/1wSBwi5wYFYmJWLiSZnNLXGjAxafY0eDBxnG8/Y4RCfQ21HvsYMe2nvNLctwY7N7sfzdv3o9d5TKbRqhF06tFM4siU6HkO47FF2FH86RPvfZRP71FBxAggw5M9w4kiegTYEz+2RwhGTByZQUEZTJSePUrMSKMkC/OW7ubm5hHN2nZ7vb5+vX79+uuvv/7682+//OMfX/7xy/98/vz555eX9dd1bZ9bsy9E61ci+kpEN/oDdv0/+iMEAET3Y5cQkfz9738vt6encimlfnp+nv7y8eNMEZeMeAr3D8H8gTM/qepHrfWnaaqfpsvl03KZPz1/eP70fHn+OD89Xeq0LFNdplK0cCm1qhYp/Z1KxKpStEp/f3oPEySPdF9yCjHLKP/twXLvGRohwtun79zI06t3x8DKe+T83Yefp4P8HgDsV/nmWP0mh0BHwPLmZ+eh5durvxkiH0eVx5t47wb2r94dR95mQc43OtoWjgDgeLz7nb97n+dHdc9wMPV+7HMAcF4F8XaA/dHz/zt+eL0+czn2FtvrtL83X8+3qdd3n8U3B8r7LZ4/H0fV/fLnFwXdV2r01SZ7ACCjo/pbcRxg722A3Gfq41aVKJNMOG2krkrPpvfv+n79mU4Z6RnhOTIBSS6RHGnpMWbpQX2A3mfzkRZhnuHhbmke1ov81CLc28j/9/l7EKWZ9cE/wsLd3foVaJQVIjPdzGgEB54Z3E/9mOEUlubhEUcNgIgoIrmPKnleNRBEyT010LMApWhRLSqiIxiovRigOiYdvUzQSwM6pvlaa48bSq37AamIiooop0jPFLAKc0qqsEhvOqicIkVZpAix9qOSyJtX5z7oj6T2EQDknjEd030V4b6raF8uH73NnVQKl31rhX3sV2VK76thuFfNJZhUlZLHar3sG/zQdwKASB9zcn6z4RL3As79RXtMBjhHOb2/uoIyOWOU8TPTkzLCg5J6rOjp5kcs2FrzzdbNttba1tzC1tY2s3VtZi3NLDxbs7bZ9npb13Zt6/pya+1LrOtni/hM7i8t81UyX5PopRK9RMSrmb3+9ttv7Xa7bT///LPRsfvT8fHPJuz+z/1RAoDv4dOHUM8WKBGVDx8+1GVZaq21Pv31r/XThw/T5XKZPvzlaS7zMs86zzxNk2ZOmTIb+SLJM6VfiORCGU9M+qQqT1rkSUu5lFKXWutSpmkptc5ay1RrrVK0Fq2lVlUtUkRKYeFyFABFmYmkbw/V03g8ovGRVJB9lRUfabU9sXdOTo8HvR/QY3TxP4TN94P+6WjPj0mDUwDw5r+8p8HfS9Px6bp5/9V+zYf+A95jnfF6P8X4b/+Lp6v1AKBXWPfU/eOKvzzt/HU/Q+DpLz3W934b5pzfdfvgx3QKco4rnC75dlXX2z/8zXN/3oQpx6/lzbv+bQAwdpx6s/xsv3Q/YB4Zo989XNwLQd8EAN+8JHJfa54S5zMO7uvt7ztVHE/LSG/3p6anZYWIKIKE+hSt193ve3WNRHtKH2xj7OGRkZHsFJHRZ/ph49fch+7w8LBIt0xn73N2C4sxjJt7c7NwM3fvI0RIjgseVYLwzDTzHjOku1kcF6AIinCPiGxu5m4R4b0UMNroer7Aws1jzO6PmJsi927SPfTJXrboW38wS/aBXkVVi4hKn1voWBvGxL0HoBRRYVWttfSagfQAYGQNSqk9BdBbCJVURUWFlUVKGdUGLkWL9m+LcI8Y5Ehh9hcjizIfOQdWEVHe0wWnfkZmFlZSojHRGafe5n4+1ZFGEO7lVU6SSN43wdnLBMKnPSnifGzY14DQMUMYXRvj5ckUPDZUDu+/HIO99f9db+2w/hLyMRNv1pqZNXdvZmZhtm1b22y7rdtqt7aur2bba7P2Ymv74q392sJekuiFgm8pcjXfbhTRiMgKkZlx29rVttbaum3t9ttv29evX7d1Xe3l5cWoRzP75/3jTzXI/8gfPQD4V+1HWqX7iqc9aKhEVGlZpo+1TpfLZZ6m5/np6TLrPM8fP36Y6zzPH5+epun5eV7meapTrXWZJladqpTKVScVmphkIaGZiSYhmYhzIaKFWGdmmUR1UtFJVGdWqaqlisiI8qWH+j3iF1WV7EH+8ffrvgQimQsxMeVYeZP3dcr70X7kJInoqMURER3df8eys/u0n8fa4qN2N9qj7ztvnYOH82z+7Sj6GAD0y7wfAOwp+MdllsdAdJ7tjj3QiYh4rIHPkRI5NnE6Xf4YdPeRafz8mGHvz0fSsVvOm3cu3x/vwyz6tGzvHIvG0evE49mM/aB3fr72NcvJtC8S3df7U+4p0+Of+V17eHDcx+n5u5dO9po9E3FQkFMSpcZIy+4nNcqkDM7e2DT2fssg3juo82gmH99kZlgSjTR9HI10sTflkR+l+sj0iMygln1Id/MI6zX6oDH6N3fziLAII08Pd29hYe4WZt4ncRHNItzJIyWVvPftx17ejySK0QSY7rHX/ZMoInrnH7m5tzBz90yP9NwDgMzsf4q7e3Lafb/hb/4hGdlTxfuSs16EF84+PVdW7ZN/4cKyr9/sg28hKlpr7w0YgUJVLcJctJR+HCi1qLKKSOGqKqx6ZBiqllq01roULaWIatG7Pl5z9PChT0iUlaXPUQqzav/V6EMYDQnMYwFkCnFfiMC96WkUEvZpDPFYAto7OY5d+mnPx2WkRZDsr6LRX9GL8j4SMRQ5YjP3CO/FfI9wD3MLD3Ozrbmt3uxm1m7ktHrEzcNfKeLazF4z6GreVvdcw7a1ma2363VdX7d1vV7Xrd3W6/V6u329vV6vn7++vLys67puRLRRX4LX6O0g/qecuf+n/H8LAP4dj9mG84dSDyQK9SbGeZqmOUuZl2VZnmq9PD8/P9VluTw9PS3L8/NluVyWp0+fLvOyLPPlMi9lmnSqtaiUOs+1aJ2K8sRSKqkWln4fnFSZpDBFIRJVosL9pPAlJIpQUSmk2UN7pdE6TOOANFYZUSYJk9BpnxoeI1CP6PdRsS9U6tdi3ceQ3g4zWg2kTwJG5/Ax5u+tFXSfKff10EdMMORRRaF9R43+NPN9F67I05X2Z30M9kQ80o/9ZzIyI3uH+V7VPN0jHUEK3V/k+/lqzne1B1L3ssvYZOqUAbnPvfd65v4H9L8v6Xz2w1P25D4TP07itAcyRONx3P+I46Ef1z6CjD7Aj61L7n8z0V6P79dlGUuiero/3VOc+z88erG0P8Kx5C5HTiB6vzyN1Po+042Isc7OvQ/nlDnK9DEm6OF9CI3Wj+QjG2vRws2aWVhztx4L9BS9uZtFho9+vtHZZ95GeiC3zYzCIszcYmQ3Co3Nl8ZKgT4L70WHoIgjxCPifX8AN/ewtPDMkYwYj42JesoiIozDI9PY72mxU/KImCicOck9iUZpZETsSdrfI5Ii43y2e38e9T0kpDAXLkWEenpeiaqo1p4pKCwiXIqUIlqlSmXW2n9QdCplKrVULbXOtc46TZOUUkspKqVoVdUczU7MLKWoVi2yTzBEtAcAPVDpxwjq66qUtTc09NF+f8VRz04R9eV4e9ZuBH0UQf0VE0T9BeKRFuEtM7eIbGHeKHJL5kbu5kxbRnqYWWQ2d2+jXNNaa81bW7dta7fr9XZbX69fX75eX19u19vLy+u6bdfX2+11/fr1er1er9Rr6yv1gdzoPjs/D+LnPYbhBxAA/Oedx5xzAMF0z0wU6hmJaXxUqnWupczzPC8islyWZZ5UF52myzxNl2VZLnWuyzzPyzRflrJMU53qvExzLdNSVKSXE6uOt3pvLhLta46VRhFQmElJSl/XKj10UC217gewftwgkmRmkpGQPFqPWUiSk1iUdNQYs2/jJCkcupfmx5FjjHNCLKzEnPvyaAq+nyOPTzWQGBN/ZiaJve3o/qyK077vfXr2eqOk9hMRK1GfvDI/vro5901Ux/30aTMf27Ds60juPR7Mcmz90Q+WeSwFpiA6zhKRct9qdT+L0/nuy5ttou4piPNlvg1i3qT4R9p+BDc9ZZNOST4GdgkiCk+jXjKljGCLsZvsPl3P0WBnaUS9Jm7u6RmeaWatD+wRzn1yZmnerDW38Gbm5m1rzWxrt21rtm3evFddzVqsa7PMbfPWcm19Gm/W0vsNuaWFu1mm8Wi2c47g4CD3YOZ0ogiOoPuAzP1t46enhFhEHrdIPNL4QZHUMw5G7uREQczB7mFEwX0wTxpJaHN3IjvtrV3O7+Mks8fZIY/L7P9gLqUo9Z3mj6KOEqmqKhGxUX/jjwUEJXsQwUREkqlSe2ugMJexNFAKc9FpqlpKnaZprlVnLaWwVhEdjQPjHa+q0uuUWoRZVbUvHRxdyazKe/tgX0A1Kpf9zXF/LNwLQpwUI0dEfbzOltas/7t7bX1bt3W73V5vt9vL7Xp9ub6+Xrdtu9q6Xrdte13X9dZau1EfsM+z8HNa/Xt19D/csrn/bxAA/HfxO58fP/af94PD3/4mf43gn376ie3Z5Kk9yeVyEb9ceJ4mmWqV2Z3NTHyaOHuhlZdloYjgqJUjgqcIjqgcNTgjuEawu0tEcK2VjZvSRoWZNSLE3dXd1ckKExcnrRzRsw6ZNQqXQlTIqZD262lSDZUixIVprI1mrtxTmyokhZRLKUWFRHkv0wtRjzlYmElYREhURFiFRFh7tpKYWbOv2tkPWvf5iworj3zGGLdZ9mLKuJyK9MYoESZRYiFVEa0qOrq2lVWLHAu2WLiUUo7Z07i/4+gpTEzj3mLkTfeHQOO8u0LEkueO7RHOjHOW33crPqdNcszUR6l0tD7HaFJP8yTO8IzszezZJ9Xm4ZnuaZ6+Z9bNbNvMzWwza2bubuu2mW3N2mZra2a0ud02b27N2xbNG4WZBbUw25q7kdnq7m2L2Mhsa2bN0jZuYSFiEtHc3dzdjdmptWBmb8zJrQURRWvNN6KgbTuqPw/vkXz4+pt0/HfeM+/dzvn2z98/Diz5zuW/53u/v79nv/3bH+tiQt++399eZp6TiGjev58mrpk6TZOM75Oozx54npNHrb2UIkTEdS/vzXPudfj9MvP4mk8/z97cfHwvIqmqx/OkqtFUo1iNrbSQ2y3XssZtq/H6+hp6vcaXL1/il19+eS+l/t4HvfMZ/ssQAPz5PQYVj1//3vc/CkYeP+TN5w8f+DmTM1PycpFLJtOy8ELEMU0yzzNXd6FloXmauPSAQ7JWriMwISKapokyk2spHKfPpRROVS79Pr55rWoEU62UmZyqnJmsmpypfPwu4vhZarKmjg7oZImQYBavtS8d7bu9KjNLYRZSVcssElFFRINcI1iYUzhGNkdSmVgiWZJDgkmJRJlZlFgyY0QN0vMNvSmUZTymvX9DeoXimPD3GVimc8bYNzb6ZJU8e907R1k+MsiDqE9kiZzCnYKNMt05zDd38s0y2NZMz9E4T30w92zN1gj3dXVxDxdxc3duLcwsGnNsrbm05uu6JhH57XbbZ2/7gJr0trZK9P0BmOg/c9D/0fHre/fz797vj67/rxxP37vsuX70o+v9O4/pn73u9wKqx99j8P4TQwAAfzTfOzD+M5f9vWDo8ev3ghuit4HO3kx6PwHA+Hqe556C7rMyzkyZiJhqlVpJKlXOTK61f6ZamYiojE7J8TOix+CGLan1mZiN9LMxB7W+eonGwbgxJ21bMHNu2xZEFCtz0O32Xir1cVa2D9b08Pl7g/R7g/l7l3n8GQAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAAA/Ff9L9Cco38U0ViFAAAAAElFTkSuQmCC"></image></svg><style>@media (prefers-color-scheme: light) { :root { filter: none; } }
@media (prefers-color-scheme: dark) { :root { filter: none; } }
</style></svg>
